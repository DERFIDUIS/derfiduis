magic
tech sky130A
magscale 1 2
timestamp 1682091667
<< error_p >>
rect -294 -264 294 298
<< nwell >>
rect -294 -264 294 298
<< pmoslvt >>
rect -200 -164 200 236
<< pdiff >>
rect -258 224 -200 236
rect -258 -152 -246 224
rect -212 -152 -200 224
rect -258 -164 -200 -152
rect 200 224 258 236
rect 200 -152 212 224
rect 246 -152 258 224
rect 200 -164 258 -152
<< pdiffc >>
rect -246 -152 -212 224
rect 212 -152 246 224
<< poly >>
rect -200 236 200 262
rect -200 -211 200 -164
rect -200 -245 -184 -211
rect 184 -245 200 -211
rect -200 -261 200 -245
<< polycont >>
rect -184 -245 184 -211
<< locali >>
rect -246 224 -212 240
rect -246 -168 -212 -152
rect 212 224 246 240
rect 212 -168 246 -152
rect -200 -245 -184 -211
rect 184 -245 200 -211
<< viali >>
rect -246 -152 -212 224
rect 212 -152 246 224
rect -184 -245 184 -211
<< metal1 >>
rect -252 224 -206 236
rect -252 -152 -246 224
rect -212 -152 -206 224
rect -252 -164 -206 -152
rect 206 224 252 236
rect 206 -152 212 224
rect 246 -152 252 224
rect 206 -164 252 -152
rect -196 -211 196 -205
rect -196 -245 -184 -211
rect 184 -245 196 -211
rect -196 -251 196 -245
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 2 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
