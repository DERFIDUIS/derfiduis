* NGSPICE file created from rectifier_lvt_01v8_end.ext - technology: sky130A

.subckt rectifier_lvt_01v8_end vinp vinn out1 vss out2
M21 a_14044_n3057# a_14114_n2960# out1 vss sky130_fd_pr__nfet_01v8_lvt ad=4.35e+12p pd=3.174e+07u as=1.8e+13p ps=1.272e+08u w=5e+06u l=180000u
M31 out2 a_14044_n3057# a_14114_n2960# out2 sky130_fd_pr__pfet_01v8_lvt ad=1.8e+13p pd=1.272e+08u as=4.35e+12p ps=3.174e+07u w=5e+06u l=350000u
M11 a_14114_n2960# a_14044_n3057# out1 vss sky130_fd_pr__nfet_01v8_lvt ad=4.35e+12p pd=3.174e+07u as=0p ps=0u w=5e+06u l=180000u
M41 a_14044_n3057# a_14114_n2960# out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=4.35e+12p pd=3.174e+07u as=0p ps=0u w=5e+06u l=350000u
M42 a_14044_n3057# a_14114_n2960# out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M22 out1 a_14114_n2960# a_14044_n3057# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M12 out1 a_14044_n3057# a_14114_n2960# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M32 a_14114_n2960# a_14044_n3057# out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M13 a_14114_n2960# a_14044_n3057# out1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M14 out1 a_14044_n3057# a_14114_n2960# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M15 a_14114_n2960# a_14044_n3057# out1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M43 out2 a_14114_n2960# a_14044_n3057# out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M33 out2 a_14044_n3057# a_14114_n2960# out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M23 a_14044_n3057# a_14114_n2960# out1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
XC2 a_14044_n3057# vinn sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
M24 out1 a_14114_n2960# a_14044_n3057# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M44 a_14044_n3057# a_14114_n2960# out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
XC1 vinp a_14114_n2960# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
XC32 out2 vss sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
M34 a_14114_n2960# a_14044_n3057# out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
XC31 out2 vss sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
M35 a_14114_n2960# a_14044_n3057# out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M16 out1 a_14044_n3057# a_14114_n2960# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M36 out2 a_14044_n3057# a_14114_n2960# out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M45 out2 a_14114_n2960# a_14044_n3057# out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M46 out2 a_14114_n2960# a_14044_n3057# out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M25 a_14044_n3057# a_14114_n2960# out1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M26 out1 a_14114_n2960# a_14044_n3057# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
.ends

