* NGSPICE file created from rectifier.ext - technology: sky130A

.subckt rectifier vinp vinn vrec vss
X0 w_13310_7310.t16 a_13470_7313.t12 a_13540_7410.t5 w_13310_7310.t15 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X1 a_730_7313.t6 a_800_7410.t13 w_n4828_7260.t26 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X2 vinp.t12 a_19910_7410.t10 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X3 a_19910_7410.t3 a_19840_7313.t12 w_13310_7310.t3 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X4 vrec.t23 a_29168_7410.t13 a_29098_7313.t11 vrec.t22 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X5 a_29098_7313.t12 vinn.t0 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X6 w_n4828_7260.t30 a_800_7410.t14 a_730_7313.t5 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X7 w_570_7310.t34 a_800_7410.t15 a_730_7313.t0 w_570_7310.t33 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X8 w_6940_7310.t19 a_13470_7313.t13 a_13540_7410.t8 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X9 w_570_7310.t17 a_730_7313.t12 a_800_7410.t6 w_570_7310.t16 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X10 w_570_7310.t32 a_800_7410.t16 a_730_7313.t7 w_570_7310.t31 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X11 a_7100_7313.t5 a_7170_7410.t13 w_6940_7310.t27 w_6940_7310.t26 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X12 vrec.t24 vss.t9 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X13 vinp.t5 vinn.t17 w_n4828_7260.t11 w_n4828_7260.t10 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X14 a_7170_7410.t8 a_7100_7313.t12 w_6940_7310.t23 w_6940_7310.t22 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X15 w_n4828_7260.t28 a_800_7410.t17 a_730_7313.t4 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X16 vinp.t1 vinn.t18 w_n4828_7260.t3 w_n4828_7260.t2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X17 vinn.t10 vinp.t13 w_n4828_7260.t35 w_n4828_7260.t34 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X18 a_730_7313.t8 a_800_7410.t18 w_570_7310.t30 w_570_7310.t29 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X19 a_800_7410.t7 a_730_7313.t13 w_570_7310.t15 w_570_7310.t14 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X20 w_6940_7310.t18 a_13470_7313.t14 a_13540_7410.t2 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X21 w_n4828_7260.t17 vinp.t14 vinn.t9 w_n4828_7260.t16 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X22 a_800_7410.t3 a_730_7313.t14 w_570_7310.t13 w_570_7310.t12 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X23 a_13470_7313.t10 a_13540_7410.t13 w_13310_7310.t35 w_13310_7310.t34 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X24 a_19840_7313.t3 a_19910_7410.t13 w_19680_7310.t17 w_19680_7310.t16 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X25 a_19910_7410.t2 a_19840_7313.t13 w_19680_7310.t29 w_19680_7310.t28 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X26 vss.t1 vinp.t15 vinn.t16 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X27 a_19840_7313.t10 a_19910_7410.t14 w_13310_7310.t1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X28 a_29098_7313.t8 a_29168_7410.t14 vrec.t21 vrec.t20 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X29 a_29168_7410.t12 a_29098_7313.t13 vrec.t11 vrec.t10 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X30 w_6940_7310.t11 a_7100_7313.t13 a_7170_7410.t4 w_6940_7310.t10 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X31 w_n4828_7260.t18 a_730_7313.t15 a_800_7410.t8 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X32 vrec.t25 vss.t8 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X33 w_13310_7310.t18 a_19910_7410.t15 a_19840_7313.t9 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X34 w_570_7310.t11 a_730_7313.t16 a_800_7410.t0 w_570_7310.t10 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X35 a_7170_7410.t10 a_7100_7313.t14 w_570_7310.t19 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X36 vss.t6 vinn.t19 vinp.t10 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X37 a_13540_7410.t4 a_13470_7313.t15 w_13310_7310.t14 w_13310_7310.t13 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X38 a_7170_7410.t3 a_7100_7313.t15 w_570_7310.t2 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X39 vss.t5 vinn.t20 vinp.t9 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X40 vrec.t9 a_29098_7313.t14 a_29168_7410.t1 vrec.t8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X41 a_19910_7410.t12 a_19840_7313.t14 w_19680_7310.t27 w_19680_7310.t26 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X42 vrec.t19 a_29168_7410.t15 a_29098_7313.t7 vrec.t18 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X43 a_7170_7410.t0 a_7100_7313.t16 w_570_7310.t1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X44 a_19910_7410.t9 a_19840_7313.t15 w_13310_7310.t21 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X45 vss.t3 vinn.t21 vinp.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X46 w_n4828_7260.t7 vinp.t16 vinn.t8 w_n4828_7260.t6 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X47 w_n4828_7260.t9 vinn.t22 vinp.t2 w_n4828_7260.t8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X48 w_13310_7310.t2 a_19840_7313.t16 a_19910_7410.t1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X49 vinp.t4 vinn.t23 vss.t2 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X50 a_730_7313.t9 a_800_7410.t19 w_570_7310.t28 w_570_7310.t27 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X51 a_29098_7313.t4 a_29168_7410.t16 w_19680_7310.t35 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X52 a_19910_7410.t7 a_19840_7313.t17 w_13310_7310.t19 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X53 a_29168_7410.t6 a_29098_7313.t15 w_19680_7310.t5 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X54 w_n4828_7260.t23 vinn.t24 vinp.t11 w_n4828_7260.t22 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X55 w_13310_7310.t33 a_13540_7410.t14 a_13470_7313.t11 w_13310_7310.t32 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X56 w_13310_7310.t12 a_13470_7313.t16 a_13540_7410.t3 w_13310_7310.t11 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X57 a_7100_7313.t11 a_7170_7410.t14 w_570_7310.t20 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X58 a_730_7313.t17 vinn.t2 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X59 w_13310_7310.t17 a_19840_7313.t18 a_19910_7410.t4 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X60 w_19680_7310.t25 a_19840_7313.t19 a_19910_7410.t5 w_19680_7310.t24 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X61 a_19840_7313.t1 a_19910_7410.t16 w_19680_7310.t15 w_19680_7310.t14 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X62 a_7100_7313.t10 a_7170_7410.t15 w_570_7310.t22 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X63 vss.t13 vinp.t17 vinn.t15 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X64 vinn.t14 vinp.t18 vss.t7 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X65 vinp.t19 a_29168_7410.t10 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X66 a_7100_7313.t9 a_7170_7410.t16 w_570_7310.t0 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X67 vss.t11 vinp.t20 vinn.t13 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X68 a_13470_7313.t17 vinn.t1 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X69 w_570_7310.t35 a_7170_7410.t17 a_7100_7313.t8 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X70 vinn.t12 vinp.t21 vss.t10 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X71 w_6940_7310.t13 a_7170_7410.t18 a_7100_7313.t4 w_6940_7310.t12 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X72 w_6940_7310.t3 a_7100_7313.t17 a_7170_7410.t2 w_6940_7310.t2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X73 w_570_7310.t26 a_800_7410.t20 a_730_7313.t11 w_570_7310.t25 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X74 a_29168_7410.t5 a_29098_7313.t16 w_19680_7310.t4 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X75 a_19840_7313.t8 a_19910_7410.t17 w_13310_7310.t20 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X76 w_570_7310.t9 a_730_7313.t18 a_800_7410.t2 w_570_7310.t8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X77 a_7170_7410.t7 a_7100_7313.t18 w_6940_7310.t21 w_6940_7310.t20 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X78 a_7100_7313.t3 a_7170_7410.t19 w_6940_7310.t7 w_6940_7310.t6 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X79 a_7100_7313.t19 vinn.t3 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X80 a_29098_7313.t6 a_29168_7410.t17 w_19680_7310.t34 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X81 w_570_7310.t5 a_7170_7410.t20 a_7100_7313.t7 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X82 vinn.t11 vinp.t22 vss.t12 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X83 a_7170_7410.t11 a_7100_7313.t20 w_6940_7310.t25 w_6940_7310.t24 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X84 vinn.t7 vinp.t23 w_n4828_7260.t15 w_n4828_7260.t14 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X85 a_19840_7313.t7 a_19910_7410.t18 w_13310_7310.t23 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X86 w_13310_7310.t22 a_19910_7410.t19 a_19840_7313.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X87 w_19680_7310.t13 a_19910_7410.t20 a_19840_7313.t2 w_19680_7310.t12 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X88 w_19680_7310.t23 a_19840_7313.t20 a_19910_7410.t8 w_19680_7310.t22 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X89 w_19680_7310.t11 a_19910_7410.t21 a_19840_7313.t0 w_19680_7310.t10 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X90 a_19840_7313.t11 a_19910_7410.t22 w_19680_7310.t9 w_19680_7310.t8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X91 w_13310_7310.t4 a_19910_7410.t23 a_19840_7313.t5 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X92 a_13470_7313.t8 a_13540_7410.t15 w_13310_7310.t31 w_13310_7310.t30 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X93 a_19910_7410.t6 a_19840_7313.t21 w_19680_7310.t21 w_19680_7310.t20 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X94 a_29168_7410.t8 a_29098_7313.t17 w_19680_7310.t3 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X95 a_29098_7313.t3 a_29168_7410.t18 vrec.t17 vrec.t16 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X96 a_29098_7313.t2 a_29168_7410.t19 w_19680_7310.t33 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X97 vinp.t7 vinn.t25 vss.t4 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X98 vrec.t7 a_29098_7313.t18 a_29168_7410.t0 vrec.t6 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X99 w_19680_7310.t32 a_29168_7410.t20 a_29098_7313.t9 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X100 w_570_7310.t4 a_7100_7313.t21 a_7170_7410.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X101 vinp.t3 vinn.t26 vss.t0 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X102 w_6940_7310.t1 a_7100_7313.t22 a_7170_7410.t1 w_6940_7310.t0 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X103 w_570_7310.t3 a_7100_7313.t23 a_7170_7410.t5 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X104 w_13310_7310.t0 a_19840_7313.t22 a_19910_7410.t0 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X105 a_800_7410.t12 a_730_7313.t19 w_n4828_7260.t25 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X106 w_13310_7310.t29 a_13540_7410.t16 a_13470_7313.t9 w_13310_7310.t28 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X107 w_19680_7310.t31 a_29168_7410.t21 a_29098_7313.t5 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X108 w_19680_7310.t2 a_29098_7313.t19 a_29168_7410.t4 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X109 a_29168_7410.t2 a_29098_7313.t20 vrec.t5 vrec.t4 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X110 a_19840_7313.t23 vinn.t4 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X111 a_29098_7313.t0 a_29168_7410.t22 vrec.t15 vrec.t14 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X112 a_7100_7313.t2 a_7170_7410.t21 w_6940_7310.t5 w_6940_7310.t4 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X113 a_29168_7410.t9 a_29098_7313.t21 vrec.t3 vrec.t2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X114 vinp.t0 vinn.t27 w_n4828_7260.t1 w_n4828_7260.t0 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X115 vinn.t6 vinp.t24 w_n4828_7260.t33 w_n4828_7260.t32 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X116 a_800_7410.t4 a_730_7313.t20 w_570_7310.t7 w_570_7310.t6 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X117 w_n4828_7260.t5 vinp.t25 vinn.t5 w_n4828_7260.t4 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X118 w_19680_7310.t1 a_29098_7313.t22 a_29168_7410.t11 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X119 a_730_7313.t3 a_800_7410.t21 w_n4828_7260.t31 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X120 w_570_7310.t21 a_7170_7410.t22 a_7100_7313.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X121 a_730_7313.t2 a_800_7410.t22 w_n4828_7260.t29 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X122 vinp.t26 a_800_7410.t10 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X123 a_13540_7410.t11 a_13470_7313.t18 w_6940_7310.t17 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X124 w_n4828_7260.t27 a_800_7410.t23 a_730_7313.t1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X125 a_13540_7410.t10 a_13470_7313.t19 w_6940_7310.t16 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X126 w_6940_7310.t15 a_13470_7313.t20 a_13540_7410.t9 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X127 vrec.t1 a_29098_7313.t23 a_29168_7410.t7 vrec.t0 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X128 w_6940_7310.t29 a_7170_7410.t23 a_7100_7313.t1 w_6940_7310.t28 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X129 w_19680_7310.t0 a_29098_7313.t24 a_29168_7410.t3 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X130 a_13540_7410.t1 a_13470_7313.t21 w_6940_7310.t14 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X131 vinp.t27 a_13540_7410.t12 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X132 w_19680_7310.t30 a_29168_7410.t23 a_29098_7313.t10 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X133 w_6940_7310.t9 a_7170_7410.t24 a_7100_7313.t0 w_6940_7310.t8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X134 vinp.t28 a_7170_7410.t12 sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X135 a_13540_7410.t0 a_13470_7313.t22 w_13310_7310.t10 w_13310_7310.t9 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X136 a_13470_7313.t4 a_13540_7410.t17 w_6940_7310.t35 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X137 w_570_7310.t18 a_7100_7313.t24 a_7170_7410.t9 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X138 w_19680_7310.t7 a_19910_7410.t24 a_19840_7313.t4 w_19680_7310.t6 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X139 a_800_7410.t9 a_730_7313.t21 w_n4828_7260.t19 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X140 vrec.t13 a_29168_7410.t24 a_29098_7313.t1 vrec.t12 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X141 w_19680_7310.t19 a_19840_7313.t24 a_19910_7410.t11 w_19680_7310.t18 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X142 a_13470_7313.t5 a_13540_7410.t18 w_6940_7310.t34 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X143 a_13540_7410.t7 a_13470_7313.t23 w_13310_7310.t8 w_13310_7310.t7 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X144 w_6940_7310.t33 a_13540_7410.t19 a_13470_7313.t0 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X145 a_13470_7313.t1 a_13540_7410.t20 w_13310_7310.t27 w_13310_7310.t26 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X146 w_n4828_7260.t13 a_730_7313.t22 a_800_7410.t5 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X147 w_6940_7310.t32 a_13540_7410.t21 a_13470_7313.t2 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X148 a_13470_7313.t3 a_13540_7410.t22 w_6940_7310.t31 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X149 a_800_7410.t1 a_730_7313.t23 w_n4828_7260.t12 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X150 a_730_7313.t10 a_800_7410.t24 w_570_7310.t24 w_570_7310.t23 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X151 w_n4828_7260.t24 a_730_7313.t24 a_800_7410.t11 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X152 w_6940_7310.t30 a_13540_7410.t23 a_13470_7313.t6 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
X153 w_n4828_7260.t21 vinn.t28 vinp.t8 w_n4828_7260.t20 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X154 w_13310_7310.t6 a_13470_7313.t24 a_13540_7410.t6 w_13310_7310.t5 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
X155 w_13310_7310.t25 a_13540_7410.t24 a_13470_7313.t7 w_13310_7310.t24 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
R0 a_13470_7313.n8 a_13470_7313.t19 708.034
R1 a_13470_7313.n7 a_13470_7313.t21 708.034
R2 a_13470_7313.n9 a_13470_7313.t18 708.034
R3 a_13470_7313.n8 a_13470_7313.t13 708.034
R4 a_13470_7313.n7 a_13470_7313.t14 708.034
R5 a_13470_7313.n9 a_13470_7313.t20 708.034
R6 a_13470_7313.n10 a_13470_7313.t23 388.664
R7 a_13470_7313.n0 a_13470_7313.t16 388.587
R8 a_13470_7313.n0 a_13470_7313.t15 388.587
R9 a_13470_7313.n6 a_13470_7313.t24 388.587
R10 a_13470_7313.n6 a_13470_7313.t22 388.587
R11 a_13470_7313.n10 a_13470_7313.t12 388.543
R12 a_13470_7313.n16 a_13470_7313.t9 5.713
R13 a_13470_7313.n16 a_13470_7313.t8 5.713
R14 a_13470_7313.n3 a_13470_7313.t7 5.713
R15 a_13470_7313.n3 a_13470_7313.t10 5.713
R16 a_13470_7313.n13 a_13470_7313.t11 5.713
R17 a_13470_7313.n13 a_13470_7313.t1 5.713
R18 a_13470_7313.n2 a_13470_7313.t2 3.48
R19 a_13470_7313.n2 a_13470_7313.t5 3.48
R20 a_13470_7313.n12 a_13470_7313.t6 3.48
R21 a_13470_7313.n12 a_13470_7313.t3 3.48
R22 a_13470_7313.t0 a_13470_7313.n18 3.48
R23 a_13470_7313.n18 a_13470_7313.t4 3.48
R24 a_13470_7313.t17 a_13470_7313.n1 2.556
R25 a_13470_7313.n1 a_13470_7313.n7 2.489
R26 a_13470_7313.n11 a_13470_7313.n9 2.478
R27 a_13470_7313.n0 a_13470_7313.n8 2.348
R28 a_13470_7313.n0 a_13470_7313.n11 0.848
R29 a_13470_7313.n1 a_13470_7313.n0 0.841
R30 a_13470_7313.n4 a_13470_7313.n2 0.701
R31 a_13470_7313.n14 a_13470_7313.n12 0.701
R32 a_13470_7313.n18 a_13470_7313.n17 0.701
R33 a_13470_7313.n14 a_13470_7313.n13 0.463
R34 a_13470_7313.n17 a_13470_7313.n16 0.463
R35 a_13470_7313.n4 a_13470_7313.n3 0.419
R36 a_13470_7313.t17 a_13470_7313.n14 0.141
R37 a_13470_7313.n15 a_13470_7313.t17 0.14
R38 a_13470_7313.n15 a_13470_7313.n5 0.135
R39 a_13470_7313.n17 a_13470_7313.n15 0.116
R40 a_13470_7313.n5 a_13470_7313.n4 0.112
R41 a_13470_7313.n11 a_13470_7313.n10 0.099
R42 a_13470_7313.n1 a_13470_7313.n6 0.077
R43 a_13540_7410.n7 a_13540_7410.t18 708.072
R44 a_13540_7410.n9 a_13540_7410.t17 708.056
R45 a_13540_7410.n11 a_13540_7410.t23 708.054
R46 a_13540_7410.n11 a_13540_7410.t22 708.054
R47 a_13540_7410.n9 a_13540_7410.t19 708.05
R48 a_13540_7410.n7 a_13540_7410.t21 708.038
R49 a_13540_7410.n6 a_13540_7410.t24 388.574
R50 a_13540_7410.n6 a_13540_7410.t13 388.524
R51 a_13540_7410.n12 a_13540_7410.t20 388.509
R52 a_13540_7410.n12 a_13540_7410.t14 388.509
R53 a_13540_7410.n10 a_13540_7410.t15 388.509
R54 a_13540_7410.n10 a_13540_7410.t16 388.509
R55 a_13540_7410.n13 a_13540_7410.t6 5.713
R56 a_13540_7410.n13 a_13540_7410.t0 5.713
R57 a_13540_7410.n5 a_13540_7410.t3 5.713
R58 a_13540_7410.n5 a_13540_7410.t4 5.713
R59 a_13540_7410.n3 a_13540_7410.t5 5.713
R60 a_13540_7410.n3 a_13540_7410.t7 5.713
R61 a_13540_7410.n4 a_13540_7410.t8 3.48
R62 a_13540_7410.n4 a_13540_7410.t10 3.48
R63 a_13540_7410.n2 a_13540_7410.t9 3.48
R64 a_13540_7410.n2 a_13540_7410.t11 3.48
R65 a_13540_7410.n14 a_13540_7410.t2 3.48
R66 a_13540_7410.t1 a_13540_7410.n14 3.48
R67 a_13540_7410.t12 a_13540_7410.n1 2.751
R68 a_13540_7410.n1 a_13540_7410.n11 2.272
R69 a_13540_7410.n8 a_13540_7410.n7 2.265
R70 a_13540_7410.n0 a_13540_7410.n9 2.178
R71 a_13540_7410.n14 a_13540_7410.n13 1.165
R72 a_13540_7410.n5 a_13540_7410.n4 1.164
R73 a_13540_7410.n3 a_13540_7410.n2 1.111
R74 a_13540_7410.n1 a_13540_7410.n0 0.841
R75 a_13540_7410.n0 a_13540_7410.n8 0.804
R76 a_13540_7410.n8 a_13540_7410.n6 0.328
R77 a_13540_7410.n1 a_13540_7410.n12 0.29
R78 a_13540_7410.t12 a_13540_7410.n3 0.2
R79 a_13540_7410.t12 a_13540_7410.n5 0.2
R80 a_13540_7410.n13 a_13540_7410.t12 0.2
R81 a_13540_7410.n0 a_13540_7410.n10 0.162
R82 w_13310_7310.n141 w_13310_7310.t24 112.822
R83 w_13310_7310.n185 w_13310_7310.t34 112.822
R84 w_13310_7310.n185 w_13310_7310.t5 112.822
R85 w_13310_7310.n261 w_13310_7310.t9 112.822
R86 w_13310_7310.n261 w_13310_7310.t28 112.822
R87 w_13310_7310.n379 w_13310_7310.t30 112.822
R88 w_13310_7310.n379 w_13310_7310.t11 112.822
R89 w_13310_7310.n455 w_13310_7310.t13 112.822
R90 w_13310_7310.n455 w_13310_7310.t32 112.822
R91 w_13310_7310.n0 w_13310_7310.t26 112.822
R92 w_13310_7310.n0 w_13310_7310.t15 112.822
R93 w_13310_7310.n45 w_13310_7310.t7 112.822
R94 w_13310_7310.n52 w_13310_7310.n49 20.699
R95 w_13310_7310.n40 w_13310_7310.n39 16.63
R96 w_13310_7310.n109 w_13310_7310.n108 16.607
R97 w_13310_7310.n423 w_13310_7310.n422 16.289
R98 w_13310_7310.n347 w_13310_7310.n346 16.289
R99 w_13310_7310.n260 w_13310_7310.n259 16.289
R100 w_13310_7310.n184 w_13310_7310.n183 16.289
R101 w_13310_7310.n500 w_13310_7310.n499 16.288
R102 w_13310_7310.n114 w_13310_7310.n110 12.641
R103 w_13310_7310.n8 w_13310_7310.n4 12.629
R104 w_13310_7310.n193 w_13310_7310.n189 12.629
R105 w_13310_7310.n269 w_13310_7310.n265 12.629
R106 w_13310_7310.n352 w_13310_7310.n348 12.629
R107 w_13310_7310.n428 w_13310_7310.n424 12.629
R108 w_13310_7310.n116 w_13310_7310.n115 9.3
R109 w_13310_7310.n122 w_13310_7310.n121 9.3
R110 w_13310_7310.n128 w_13310_7310.n127 9.3
R111 w_13310_7310.n134 w_13310_7310.n133 9.3
R112 w_13310_7310.n140 w_13310_7310.n139 9.3
R113 w_13310_7310.n152 w_13310_7310.n151 9.3
R114 w_13310_7310.n158 w_13310_7310.n157 9.3
R115 w_13310_7310.n164 w_13310_7310.n163 9.3
R116 w_13310_7310.n170 w_13310_7310.n169 9.3
R117 w_13310_7310.n176 w_13310_7310.n175 9.3
R118 w_13310_7310.n181 w_13310_7310.n180 9.3
R119 w_13310_7310.n195 w_13310_7310.n194 9.3
R120 w_13310_7310.n201 w_13310_7310.n200 9.3
R121 w_13310_7310.n207 w_13310_7310.n206 9.3
R122 w_13310_7310.n213 w_13310_7310.n212 9.3
R123 w_13310_7310.n219 w_13310_7310.n218 9.3
R124 w_13310_7310.n227 w_13310_7310.n226 9.3
R125 w_13310_7310.n233 w_13310_7310.n232 9.3
R126 w_13310_7310.n239 w_13310_7310.n238 9.3
R127 w_13310_7310.n245 w_13310_7310.n244 9.3
R128 w_13310_7310.n251 w_13310_7310.n250 9.3
R129 w_13310_7310.n256 w_13310_7310.n255 9.3
R130 w_13310_7310.n271 w_13310_7310.n270 9.3
R131 w_13310_7310.n277 w_13310_7310.n276 9.3
R132 w_13310_7310.n283 w_13310_7310.n282 9.3
R133 w_13310_7310.n289 w_13310_7310.n288 9.3
R134 w_13310_7310.n295 w_13310_7310.n294 9.3
R135 w_13310_7310.n303 w_13310_7310.n302 9.3
R136 w_13310_7310.n309 w_13310_7310.n308 9.3
R137 w_13310_7310.n315 w_13310_7310.n314 9.3
R138 w_13310_7310.n321 w_13310_7310.n320 9.3
R139 w_13310_7310.n327 w_13310_7310.n326 9.3
R140 w_13310_7310.n332 w_13310_7310.n331 9.3
R141 w_13310_7310.n354 w_13310_7310.n353 9.3
R142 w_13310_7310.n360 w_13310_7310.n359 9.3
R143 w_13310_7310.n366 w_13310_7310.n365 9.3
R144 w_13310_7310.n372 w_13310_7310.n371 9.3
R145 w_13310_7310.n378 w_13310_7310.n377 9.3
R146 w_13310_7310.n390 w_13310_7310.n389 9.3
R147 w_13310_7310.n396 w_13310_7310.n395 9.3
R148 w_13310_7310.n402 w_13310_7310.n401 9.3
R149 w_13310_7310.n408 w_13310_7310.n407 9.3
R150 w_13310_7310.n414 w_13310_7310.n413 9.3
R151 w_13310_7310.n419 w_13310_7310.n418 9.3
R152 w_13310_7310.n430 w_13310_7310.n429 9.3
R153 w_13310_7310.n436 w_13310_7310.n435 9.3
R154 w_13310_7310.n442 w_13310_7310.n441 9.3
R155 w_13310_7310.n448 w_13310_7310.n447 9.3
R156 w_13310_7310.n454 w_13310_7310.n453 9.3
R157 w_13310_7310.n466 w_13310_7310.n465 9.3
R158 w_13310_7310.n472 w_13310_7310.n471 9.3
R159 w_13310_7310.n478 w_13310_7310.n477 9.3
R160 w_13310_7310.n484 w_13310_7310.n483 9.3
R161 w_13310_7310.n490 w_13310_7310.n489 9.3
R162 w_13310_7310.n495 w_13310_7310.n494 9.3
R163 w_13310_7310.n434 w_13310_7310.n433 9.3
R164 w_13310_7310.n440 w_13310_7310.n439 9.3
R165 w_13310_7310.n446 w_13310_7310.n445 9.3
R166 w_13310_7310.n452 w_13310_7310.n451 9.3
R167 w_13310_7310.n470 w_13310_7310.n469 9.3
R168 w_13310_7310.n476 w_13310_7310.n475 9.3
R169 w_13310_7310.n482 w_13310_7310.n481 9.3
R170 w_13310_7310.n488 w_13310_7310.n487 9.3
R171 w_13310_7310.n493 w_13310_7310.n492 9.3
R172 w_13310_7310.n358 w_13310_7310.n357 9.3
R173 w_13310_7310.n364 w_13310_7310.n363 9.3
R174 w_13310_7310.n370 w_13310_7310.n369 9.3
R175 w_13310_7310.n376 w_13310_7310.n375 9.3
R176 w_13310_7310.n394 w_13310_7310.n393 9.3
R177 w_13310_7310.n400 w_13310_7310.n399 9.3
R178 w_13310_7310.n406 w_13310_7310.n405 9.3
R179 w_13310_7310.n412 w_13310_7310.n411 9.3
R180 w_13310_7310.n417 w_13310_7310.n416 9.3
R181 w_13310_7310.n275 w_13310_7310.n274 9.3
R182 w_13310_7310.n281 w_13310_7310.n280 9.3
R183 w_13310_7310.n287 w_13310_7310.n286 9.3
R184 w_13310_7310.n293 w_13310_7310.n292 9.3
R185 w_13310_7310.n307 w_13310_7310.n306 9.3
R186 w_13310_7310.n313 w_13310_7310.n312 9.3
R187 w_13310_7310.n319 w_13310_7310.n318 9.3
R188 w_13310_7310.n325 w_13310_7310.n324 9.3
R189 w_13310_7310.n330 w_13310_7310.n329 9.3
R190 w_13310_7310.n199 w_13310_7310.n198 9.3
R191 w_13310_7310.n205 w_13310_7310.n204 9.3
R192 w_13310_7310.n211 w_13310_7310.n210 9.3
R193 w_13310_7310.n217 w_13310_7310.n216 9.3
R194 w_13310_7310.n231 w_13310_7310.n230 9.3
R195 w_13310_7310.n237 w_13310_7310.n236 9.3
R196 w_13310_7310.n243 w_13310_7310.n242 9.3
R197 w_13310_7310.n249 w_13310_7310.n248 9.3
R198 w_13310_7310.n254 w_13310_7310.n253 9.3
R199 w_13310_7310.n120 w_13310_7310.n119 9.3
R200 w_13310_7310.n126 w_13310_7310.n125 9.3
R201 w_13310_7310.n132 w_13310_7310.n131 9.3
R202 w_13310_7310.n138 w_13310_7310.n137 9.3
R203 w_13310_7310.n156 w_13310_7310.n155 9.3
R204 w_13310_7310.n162 w_13310_7310.n161 9.3
R205 w_13310_7310.n168 w_13310_7310.n167 9.3
R206 w_13310_7310.n174 w_13310_7310.n173 9.3
R207 w_13310_7310.n179 w_13310_7310.n178 9.3
R208 w_13310_7310.n106 w_13310_7310.n105 9.3
R209 w_13310_7310.n54 w_13310_7310.n53 9.3
R210 w_13310_7310.n57 w_13310_7310.n56 9.3
R211 w_13310_7310.n59 w_13310_7310.n58 9.3
R212 w_13310_7310.n62 w_13310_7310.n61 9.3
R213 w_13310_7310.n64 w_13310_7310.n63 9.3
R214 w_13310_7310.n67 w_13310_7310.n66 9.3
R215 w_13310_7310.n69 w_13310_7310.n68 9.3
R216 w_13310_7310.n72 w_13310_7310.n71 9.3
R217 w_13310_7310.n74 w_13310_7310.n73 9.3
R218 w_13310_7310.n81 w_13310_7310.n80 9.3
R219 w_13310_7310.n84 w_13310_7310.n83 9.3
R220 w_13310_7310.n86 w_13310_7310.n85 9.3
R221 w_13310_7310.n89 w_13310_7310.n88 9.3
R222 w_13310_7310.n91 w_13310_7310.n90 9.3
R223 w_13310_7310.n94 w_13310_7310.n93 9.3
R224 w_13310_7310.n96 w_13310_7310.n95 9.3
R225 w_13310_7310.n99 w_13310_7310.n98 9.3
R226 w_13310_7310.n101 w_13310_7310.n100 9.3
R227 w_13310_7310.n104 w_13310_7310.n103 9.3
R228 w_13310_7310.n10 w_13310_7310.n9 9.3
R229 w_13310_7310.n14 w_13310_7310.n13 9.3
R230 w_13310_7310.n16 w_13310_7310.n15 9.3
R231 w_13310_7310.n20 w_13310_7310.n19 9.3
R232 w_13310_7310.n22 w_13310_7310.n21 9.3
R233 w_13310_7310.n26 w_13310_7310.n25 9.3
R234 w_13310_7310.n28 w_13310_7310.n27 9.3
R235 w_13310_7310.n32 w_13310_7310.n31 9.3
R236 w_13310_7310.n34 w_13310_7310.n33 9.3
R237 w_13310_7310.n532 w_13310_7310.n531 9.3
R238 w_13310_7310.n530 w_13310_7310.n529 9.3
R239 w_13310_7310.n526 w_13310_7310.n525 9.3
R240 w_13310_7310.n524 w_13310_7310.n523 9.3
R241 w_13310_7310.n520 w_13310_7310.n519 9.3
R242 w_13310_7310.n518 w_13310_7310.n517 9.3
R243 w_13310_7310.n514 w_13310_7310.n513 9.3
R244 w_13310_7310.n512 w_13310_7310.n511 9.3
R245 w_13310_7310.n508 w_13310_7310.n507 9.3
R246 w_13310_7310.n506 w_13310_7310.n505 9.3
R247 w_13310_7310.n503 w_13310_7310.n502 9.3
R248 w_13310_7310.n7 w_13310_7310.n6 8.855
R249 w_13310_7310.n427 w_13310_7310.n426 8.855
R250 w_13310_7310.n433 w_13310_7310.n432 8.855
R251 w_13310_7310.n439 w_13310_7310.n438 8.855
R252 w_13310_7310.n445 w_13310_7310.n444 8.855
R253 w_13310_7310.n451 w_13310_7310.n450 8.855
R254 w_13310_7310.n458 w_13310_7310.n457 8.855
R255 w_13310_7310.n463 w_13310_7310.n462 8.855
R256 w_13310_7310.n469 w_13310_7310.n468 8.855
R257 w_13310_7310.n475 w_13310_7310.n474 8.855
R258 w_13310_7310.n481 w_13310_7310.n480 8.855
R259 w_13310_7310.n487 w_13310_7310.n486 8.855
R260 w_13310_7310.n492 w_13310_7310.n491 8.855
R261 w_13310_7310.n351 w_13310_7310.n350 8.855
R262 w_13310_7310.n357 w_13310_7310.n356 8.855
R263 w_13310_7310.n363 w_13310_7310.n362 8.855
R264 w_13310_7310.n369 w_13310_7310.n368 8.855
R265 w_13310_7310.n375 w_13310_7310.n374 8.855
R266 w_13310_7310.n382 w_13310_7310.n381 8.855
R267 w_13310_7310.n387 w_13310_7310.n386 8.855
R268 w_13310_7310.n393 w_13310_7310.n392 8.855
R269 w_13310_7310.n399 w_13310_7310.n398 8.855
R270 w_13310_7310.n405 w_13310_7310.n404 8.855
R271 w_13310_7310.n411 w_13310_7310.n410 8.855
R272 w_13310_7310.n416 w_13310_7310.n415 8.855
R273 w_13310_7310.n268 w_13310_7310.n267 8.855
R274 w_13310_7310.n274 w_13310_7310.n273 8.855
R275 w_13310_7310.n280 w_13310_7310.n279 8.855
R276 w_13310_7310.n286 w_13310_7310.n285 8.855
R277 w_13310_7310.n292 w_13310_7310.n291 8.855
R278 w_13310_7310.n264 w_13310_7310.n263 8.855
R279 w_13310_7310.n300 w_13310_7310.n299 8.855
R280 w_13310_7310.n306 w_13310_7310.n305 8.855
R281 w_13310_7310.n312 w_13310_7310.n311 8.855
R282 w_13310_7310.n318 w_13310_7310.n317 8.855
R283 w_13310_7310.n324 w_13310_7310.n323 8.855
R284 w_13310_7310.n329 w_13310_7310.n328 8.855
R285 w_13310_7310.n192 w_13310_7310.n191 8.855
R286 w_13310_7310.n198 w_13310_7310.n197 8.855
R287 w_13310_7310.n204 w_13310_7310.n203 8.855
R288 w_13310_7310.n210 w_13310_7310.n209 8.855
R289 w_13310_7310.n216 w_13310_7310.n215 8.855
R290 w_13310_7310.n188 w_13310_7310.n187 8.855
R291 w_13310_7310.n224 w_13310_7310.n223 8.855
R292 w_13310_7310.n230 w_13310_7310.n229 8.855
R293 w_13310_7310.n236 w_13310_7310.n235 8.855
R294 w_13310_7310.n242 w_13310_7310.n241 8.855
R295 w_13310_7310.n248 w_13310_7310.n247 8.855
R296 w_13310_7310.n253 w_13310_7310.n252 8.855
R297 w_13310_7310.n113 w_13310_7310.n112 8.855
R298 w_13310_7310.n119 w_13310_7310.n118 8.855
R299 w_13310_7310.n125 w_13310_7310.n124 8.855
R300 w_13310_7310.n131 w_13310_7310.n130 8.855
R301 w_13310_7310.n137 w_13310_7310.n136 8.855
R302 w_13310_7310.n144 w_13310_7310.n143 8.855
R303 w_13310_7310.n149 w_13310_7310.n148 8.855
R304 w_13310_7310.n155 w_13310_7310.n154 8.855
R305 w_13310_7310.n161 w_13310_7310.n160 8.855
R306 w_13310_7310.n167 w_13310_7310.n166 8.855
R307 w_13310_7310.n173 w_13310_7310.n172 8.855
R308 w_13310_7310.n178 w_13310_7310.n177 8.855
R309 w_13310_7310.n51 w_13310_7310.n50 8.855
R310 w_13310_7310.n56 w_13310_7310.n55 8.855
R311 w_13310_7310.n61 w_13310_7310.n60 8.855
R312 w_13310_7310.n66 w_13310_7310.n65 8.855
R313 w_13310_7310.n71 w_13310_7310.n70 8.855
R314 w_13310_7310.n76 w_13310_7310.n75 8.855
R315 w_13310_7310.n48 w_13310_7310.n47 8.855
R316 w_13310_7310.n83 w_13310_7310.n82 8.855
R317 w_13310_7310.n88 w_13310_7310.n87 8.855
R318 w_13310_7310.n93 w_13310_7310.n92 8.855
R319 w_13310_7310.n98 w_13310_7310.n97 8.855
R320 w_13310_7310.n103 w_13310_7310.n102 8.855
R321 w_13310_7310.n13 w_13310_7310.n12 8.855
R322 w_13310_7310.n19 w_13310_7310.n18 8.855
R323 w_13310_7310.n25 w_13310_7310.n24 8.855
R324 w_13310_7310.n31 w_13310_7310.n30 8.855
R325 w_13310_7310.n3 w_13310_7310.n2 8.855
R326 w_13310_7310.n38 w_13310_7310.n37 8.855
R327 w_13310_7310.n529 w_13310_7310.n528 8.855
R328 w_13310_7310.n523 w_13310_7310.n522 8.855
R329 w_13310_7310.n517 w_13310_7310.n516 8.855
R330 w_13310_7310.n511 w_13310_7310.n510 8.855
R331 w_13310_7310.n505 w_13310_7310.n504 8.855
R332 w_13310_7310.n47 w_13310_7310.n46 7.775
R333 w_13310_7310.n496 w_13310_7310.n423 6.209
R334 w_13310_7310.n420 w_13310_7310.n347 6.209
R335 w_13310_7310.n333 w_13310_7310.n260 6.209
R336 w_13310_7310.n257 w_13310_7310.n184 6.209
R337 w_13310_7310.n501 w_13310_7310.n500 6.209
R338 w_13310_7310.n182 w_13310_7310.n109 6.208
R339 w_13310_7310.n456 w_13310_7310.n455 5.95
R340 w_13310_7310.n380 w_13310_7310.n379 5.95
R341 w_13310_7310.n262 w_13310_7310.n261 5.95
R342 w_13310_7310.n186 w_13310_7310.n185 5.95
R343 w_13310_7310.n1 w_13310_7310.n0 5.95
R344 w_13310_7310.n464 w_13310_7310.n463 5.876
R345 w_13310_7310.n388 w_13310_7310.n387 5.876
R346 w_13310_7310.n301 w_13310_7310.n300 5.876
R347 w_13310_7310.n225 w_13310_7310.n224 5.876
R348 w_13310_7310.n533 w_13310_7310.n38 5.876
R349 w_13310_7310.n77 w_13310_7310.n76 5.873
R350 w_13310_7310.n150 w_13310_7310.n149 5.873
R351 w_13310_7310.n534 w_13310_7310.t27 5.713
R352 w_13310_7310.n78 w_13310_7310.t8 5.713
R353 w_13310_7310.n384 w_13310_7310.t31 5.713
R354 w_13310_7310.n384 w_13310_7310.t12 5.713
R355 w_13310_7310.n146 w_13310_7310.t25 5.713
R356 w_13310_7310.n221 w_13310_7310.t35 5.713
R357 w_13310_7310.n221 w_13310_7310.t6 5.713
R358 w_13310_7310.n297 w_13310_7310.t10 5.713
R359 w_13310_7310.n297 w_13310_7310.t29 5.713
R360 w_13310_7310.n460 w_13310_7310.t14 5.713
R361 w_13310_7310.n460 w_13310_7310.t33 5.713
R362 w_13310_7310.t16 w_13310_7310.n534 5.713
R363 w_13310_7310.n107 w_13310_7310.n40 5.637
R364 w_13310_7310.n193 w_13310_7310.n192 5.614
R365 w_13310_7310.n269 w_13310_7310.n268 5.614
R366 w_13310_7310.n428 w_13310_7310.n427 5.614
R367 w_13310_7310.n352 w_13310_7310.n351 5.614
R368 w_13310_7310.n8 w_13310_7310.n7 5.614
R369 w_13310_7310.n114 w_13310_7310.n113 5.611
R370 w_13310_7310.n52 w_13310_7310.n51 5.571
R371 w_13310_7310.n142 w_13310_7310.n141 5.347
R372 w_13310_7310.n335 w_13310_7310.t18 4.491
R373 w_13310_7310.n335 w_13310_7310.t1 4.386
R374 w_13310_7310.n336 w_13310_7310.t0 4.386
R375 w_13310_7310.n337 w_13310_7310.t21 4.386
R376 w_13310_7310.n338 w_13310_7310.t4 4.386
R377 w_13310_7310.n339 w_13310_7310.t23 4.386
R378 w_13310_7310.n340 w_13310_7310.t2 4.386
R379 w_13310_7310.n341 w_13310_7310.t3 4.386
R380 w_13310_7310.n342 w_13310_7310.t22 4.386
R381 w_13310_7310.n343 w_13310_7310.t20 4.386
R382 w_13310_7310.n344 w_13310_7310.t17 4.386
R383 w_13310_7310.n345 w_13310_7310.t19 4.386
R384 w_13310_7310.n383 w_13310_7310.n382 4.27
R385 w_13310_7310.n459 w_13310_7310.n458 4.27
R386 w_13310_7310.n296 w_13310_7310.n264 4.27
R387 w_13310_7310.n220 w_13310_7310.n188 4.27
R388 w_13310_7310.n35 w_13310_7310.n3 4.27
R389 w_13310_7310.n145 w_13310_7310.n144 4.269
R390 w_13310_7310.n79 w_13310_7310.n48 4.269
R391 w_13310_7310.n172 w_13310_7310.n171 3.685
R392 w_13310_7310.n166 w_13310_7310.n165 3.685
R393 w_13310_7310.n160 w_13310_7310.n159 3.685
R394 w_13310_7310.n154 w_13310_7310.n153 3.685
R395 w_13310_7310.n148 w_13310_7310.n147 3.685
R396 w_13310_7310.n143 w_13310_7310.n142 3.685
R397 w_13310_7310.n136 w_13310_7310.n135 3.685
R398 w_13310_7310.n130 w_13310_7310.n129 3.685
R399 w_13310_7310.n124 w_13310_7310.n123 3.685
R400 w_13310_7310.n118 w_13310_7310.n117 3.685
R401 w_13310_7310.n112 w_13310_7310.n111 3.514
R402 w_13310_7310.n247 w_13310_7310.n246 3.052
R403 w_13310_7310.n241 w_13310_7310.n240 3.052
R404 w_13310_7310.n235 w_13310_7310.n234 3.052
R405 w_13310_7310.n229 w_13310_7310.n228 3.052
R406 w_13310_7310.n223 w_13310_7310.n222 3.052
R407 w_13310_7310.n187 w_13310_7310.n186 3.052
R408 w_13310_7310.n215 w_13310_7310.n214 3.052
R409 w_13310_7310.n209 w_13310_7310.n208 3.052
R410 w_13310_7310.n203 w_13310_7310.n202 3.052
R411 w_13310_7310.n197 w_13310_7310.n196 3.052
R412 w_13310_7310.n323 w_13310_7310.n322 3.052
R413 w_13310_7310.n317 w_13310_7310.n316 3.052
R414 w_13310_7310.n311 w_13310_7310.n310 3.052
R415 w_13310_7310.n305 w_13310_7310.n304 3.052
R416 w_13310_7310.n299 w_13310_7310.n298 3.052
R417 w_13310_7310.n263 w_13310_7310.n262 3.052
R418 w_13310_7310.n291 w_13310_7310.n290 3.052
R419 w_13310_7310.n285 w_13310_7310.n284 3.052
R420 w_13310_7310.n279 w_13310_7310.n278 3.052
R421 w_13310_7310.n273 w_13310_7310.n272 3.052
R422 w_13310_7310.n410 w_13310_7310.n409 3.052
R423 w_13310_7310.n404 w_13310_7310.n403 3.052
R424 w_13310_7310.n398 w_13310_7310.n397 3.052
R425 w_13310_7310.n392 w_13310_7310.n391 3.052
R426 w_13310_7310.n386 w_13310_7310.n385 3.052
R427 w_13310_7310.n381 w_13310_7310.n380 3.052
R428 w_13310_7310.n374 w_13310_7310.n373 3.052
R429 w_13310_7310.n368 w_13310_7310.n367 3.052
R430 w_13310_7310.n362 w_13310_7310.n361 3.052
R431 w_13310_7310.n356 w_13310_7310.n355 3.052
R432 w_13310_7310.n486 w_13310_7310.n485 3.052
R433 w_13310_7310.n480 w_13310_7310.n479 3.052
R434 w_13310_7310.n474 w_13310_7310.n473 3.052
R435 w_13310_7310.n468 w_13310_7310.n467 3.052
R436 w_13310_7310.n462 w_13310_7310.n461 3.052
R437 w_13310_7310.n457 w_13310_7310.n456 3.052
R438 w_13310_7310.n450 w_13310_7310.n449 3.052
R439 w_13310_7310.n444 w_13310_7310.n443 3.052
R440 w_13310_7310.n438 w_13310_7310.n437 3.052
R441 w_13310_7310.n432 w_13310_7310.n431 3.052
R442 w_13310_7310.n510 w_13310_7310.n509 3.052
R443 w_13310_7310.n516 w_13310_7310.n515 3.052
R444 w_13310_7310.n522 w_13310_7310.n521 3.052
R445 w_13310_7310.n528 w_13310_7310.n527 3.052
R446 w_13310_7310.n37 w_13310_7310.n36 3.052
R447 w_13310_7310.n2 w_13310_7310.n1 3.052
R448 w_13310_7310.n30 w_13310_7310.n29 3.052
R449 w_13310_7310.n24 w_13310_7310.n23 3.052
R450 w_13310_7310.n18 w_13310_7310.n17 3.052
R451 w_13310_7310.n12 w_13310_7310.n11 3.052
R452 w_13310_7310.n191 w_13310_7310.n190 2.91
R453 w_13310_7310.n267 w_13310_7310.n266 2.91
R454 w_13310_7310.n350 w_13310_7310.n349 2.91
R455 w_13310_7310.n426 w_13310_7310.n425 2.91
R456 w_13310_7310.n6 w_13310_7310.n5 2.91
R457 w_13310_7310.n421 w_13310_7310.n345 2.351
R458 w_13310_7310.n498 w_13310_7310.n107 0.768
R459 w_13310_7310.n258 w_13310_7310.n182 0.75
R460 w_13310_7310.n54 w_13310_7310.n52 0.713
R461 w_13310_7310.n116 w_13310_7310.n114 0.668
R462 w_13310_7310.n10 w_13310_7310.n8 0.652
R463 w_13310_7310.n195 w_13310_7310.n193 0.652
R464 w_13310_7310.n271 w_13310_7310.n269 0.652
R465 w_13310_7310.n354 w_13310_7310.n352 0.652
R466 w_13310_7310.n430 w_13310_7310.n428 0.652
R467 w_13310_7310.n334 w_13310_7310.n258 0.57
R468 w_13310_7310.n497 w_13310_7310.n421 0.57
R469 w_13310_7310.n421 w_13310_7310.n334 0.57
R470 w_13310_7310.n498 w_13310_7310.n497 0.57
R471 w_13310_7310.n45 w_13310_7310.n44 0.54
R472 w_13310_7310.n45 w_13310_7310.n43 0.54
R473 w_13310_7310.n46 w_13310_7310.n45 0.54
R474 w_13310_7310.n45 w_13310_7310.n42 0.54
R475 w_13310_7310.n45 w_13310_7310.n41 0.54
R476 w_13310_7310.n258 w_13310_7310.n257 0.208
R477 w_13310_7310.n334 w_13310_7310.n333 0.208
R478 w_13310_7310.n421 w_13310_7310.n420 0.208
R479 w_13310_7310.n497 w_13310_7310.n496 0.208
R480 w_13310_7310.n501 w_13310_7310.n498 0.208
R481 w_13310_7310.n337 w_13310_7310.n336 0.106
R482 w_13310_7310.n339 w_13310_7310.n338 0.106
R483 w_13310_7310.n341 w_13310_7310.n340 0.106
R484 w_13310_7310.n343 w_13310_7310.n342 0.106
R485 w_13310_7310.n345 w_13310_7310.n344 0.106
R486 w_13310_7310.n336 w_13310_7310.n335 0.083
R487 w_13310_7310.n338 w_13310_7310.n337 0.083
R488 w_13310_7310.n340 w_13310_7310.n339 0.083
R489 w_13310_7310.n342 w_13310_7310.n341 0.083
R490 w_13310_7310.n344 w_13310_7310.n343 0.083
R491 w_13310_7310.n152 w_13310_7310.n150 0.047
R492 w_13310_7310.n77 w_13310_7310.n74 0.046
R493 w_13310_7310.n107 w_13310_7310.n106 0.045
R494 w_13310_7310.n145 w_13310_7310.n140 0.043
R495 w_13310_7310.n81 w_13310_7310.n79 0.042
R496 w_13310_7310.n182 w_13310_7310.n181 0.04
R497 w_13310_7310.n181 w_13310_7310.n179 0.032
R498 w_13310_7310.n179 w_13310_7310.n176 0.032
R499 w_13310_7310.n176 w_13310_7310.n174 0.032
R500 w_13310_7310.n174 w_13310_7310.n170 0.032
R501 w_13310_7310.n170 w_13310_7310.n168 0.032
R502 w_13310_7310.n168 w_13310_7310.n164 0.032
R503 w_13310_7310.n164 w_13310_7310.n162 0.032
R504 w_13310_7310.n162 w_13310_7310.n158 0.032
R505 w_13310_7310.n158 w_13310_7310.n156 0.032
R506 w_13310_7310.n156 w_13310_7310.n152 0.032
R507 w_13310_7310.n140 w_13310_7310.n138 0.032
R508 w_13310_7310.n138 w_13310_7310.n134 0.032
R509 w_13310_7310.n134 w_13310_7310.n132 0.032
R510 w_13310_7310.n132 w_13310_7310.n128 0.032
R511 w_13310_7310.n128 w_13310_7310.n126 0.032
R512 w_13310_7310.n126 w_13310_7310.n122 0.032
R513 w_13310_7310.n122 w_13310_7310.n120 0.032
R514 w_13310_7310.n120 w_13310_7310.n116 0.032
R515 w_13310_7310.n227 w_13310_7310.n225 0.031
R516 w_13310_7310.n303 w_13310_7310.n301 0.031
R517 w_13310_7310.n390 w_13310_7310.n388 0.031
R518 w_13310_7310.n466 w_13310_7310.n464 0.031
R519 w_13310_7310.n533 w_13310_7310.n532 0.031
R520 w_13310_7310.n106 w_13310_7310.n104 0.031
R521 w_13310_7310.n104 w_13310_7310.n101 0.031
R522 w_13310_7310.n101 w_13310_7310.n99 0.031
R523 w_13310_7310.n99 w_13310_7310.n96 0.031
R524 w_13310_7310.n96 w_13310_7310.n94 0.031
R525 w_13310_7310.n94 w_13310_7310.n91 0.031
R526 w_13310_7310.n91 w_13310_7310.n89 0.031
R527 w_13310_7310.n89 w_13310_7310.n86 0.031
R528 w_13310_7310.n86 w_13310_7310.n84 0.031
R529 w_13310_7310.n84 w_13310_7310.n81 0.031
R530 w_13310_7310.n74 w_13310_7310.n72 0.031
R531 w_13310_7310.n72 w_13310_7310.n69 0.031
R532 w_13310_7310.n69 w_13310_7310.n67 0.031
R533 w_13310_7310.n67 w_13310_7310.n64 0.031
R534 w_13310_7310.n64 w_13310_7310.n62 0.031
R535 w_13310_7310.n62 w_13310_7310.n59 0.031
R536 w_13310_7310.n59 w_13310_7310.n57 0.031
R537 w_13310_7310.n57 w_13310_7310.n54 0.031
R538 w_13310_7310.n150 w_13310_7310.n146 0.031
R539 w_13310_7310.n78 w_13310_7310.n77 0.03
R540 w_13310_7310.n220 w_13310_7310.n219 0.029
R541 w_13310_7310.n296 w_13310_7310.n295 0.029
R542 w_13310_7310.n383 w_13310_7310.n378 0.029
R543 w_13310_7310.n459 w_13310_7310.n454 0.029
R544 w_13310_7310.n35 w_13310_7310.n34 0.029
R545 w_13310_7310.n257 w_13310_7310.n256 0.027
R546 w_13310_7310.n333 w_13310_7310.n332 0.027
R547 w_13310_7310.n420 w_13310_7310.n419 0.027
R548 w_13310_7310.n496 w_13310_7310.n495 0.027
R549 w_13310_7310.n503 w_13310_7310.n501 0.027
R550 w_13310_7310.n256 w_13310_7310.n254 0.021
R551 w_13310_7310.n254 w_13310_7310.n251 0.021
R552 w_13310_7310.n251 w_13310_7310.n249 0.021
R553 w_13310_7310.n249 w_13310_7310.n245 0.021
R554 w_13310_7310.n245 w_13310_7310.n243 0.021
R555 w_13310_7310.n243 w_13310_7310.n239 0.021
R556 w_13310_7310.n239 w_13310_7310.n237 0.021
R557 w_13310_7310.n237 w_13310_7310.n233 0.021
R558 w_13310_7310.n233 w_13310_7310.n231 0.021
R559 w_13310_7310.n231 w_13310_7310.n227 0.021
R560 w_13310_7310.n219 w_13310_7310.n217 0.021
R561 w_13310_7310.n217 w_13310_7310.n213 0.021
R562 w_13310_7310.n213 w_13310_7310.n211 0.021
R563 w_13310_7310.n211 w_13310_7310.n207 0.021
R564 w_13310_7310.n207 w_13310_7310.n205 0.021
R565 w_13310_7310.n205 w_13310_7310.n201 0.021
R566 w_13310_7310.n201 w_13310_7310.n199 0.021
R567 w_13310_7310.n199 w_13310_7310.n195 0.021
R568 w_13310_7310.n332 w_13310_7310.n330 0.021
R569 w_13310_7310.n330 w_13310_7310.n327 0.021
R570 w_13310_7310.n327 w_13310_7310.n325 0.021
R571 w_13310_7310.n325 w_13310_7310.n321 0.021
R572 w_13310_7310.n321 w_13310_7310.n319 0.021
R573 w_13310_7310.n319 w_13310_7310.n315 0.021
R574 w_13310_7310.n315 w_13310_7310.n313 0.021
R575 w_13310_7310.n313 w_13310_7310.n309 0.021
R576 w_13310_7310.n309 w_13310_7310.n307 0.021
R577 w_13310_7310.n307 w_13310_7310.n303 0.021
R578 w_13310_7310.n295 w_13310_7310.n293 0.021
R579 w_13310_7310.n293 w_13310_7310.n289 0.021
R580 w_13310_7310.n289 w_13310_7310.n287 0.021
R581 w_13310_7310.n287 w_13310_7310.n283 0.021
R582 w_13310_7310.n283 w_13310_7310.n281 0.021
R583 w_13310_7310.n281 w_13310_7310.n277 0.021
R584 w_13310_7310.n277 w_13310_7310.n275 0.021
R585 w_13310_7310.n275 w_13310_7310.n271 0.021
R586 w_13310_7310.n419 w_13310_7310.n417 0.021
R587 w_13310_7310.n417 w_13310_7310.n414 0.021
R588 w_13310_7310.n414 w_13310_7310.n412 0.021
R589 w_13310_7310.n412 w_13310_7310.n408 0.021
R590 w_13310_7310.n408 w_13310_7310.n406 0.021
R591 w_13310_7310.n406 w_13310_7310.n402 0.021
R592 w_13310_7310.n402 w_13310_7310.n400 0.021
R593 w_13310_7310.n400 w_13310_7310.n396 0.021
R594 w_13310_7310.n396 w_13310_7310.n394 0.021
R595 w_13310_7310.n394 w_13310_7310.n390 0.021
R596 w_13310_7310.n378 w_13310_7310.n376 0.021
R597 w_13310_7310.n376 w_13310_7310.n372 0.021
R598 w_13310_7310.n372 w_13310_7310.n370 0.021
R599 w_13310_7310.n370 w_13310_7310.n366 0.021
R600 w_13310_7310.n366 w_13310_7310.n364 0.021
R601 w_13310_7310.n364 w_13310_7310.n360 0.021
R602 w_13310_7310.n360 w_13310_7310.n358 0.021
R603 w_13310_7310.n358 w_13310_7310.n354 0.021
R604 w_13310_7310.n495 w_13310_7310.n493 0.021
R605 w_13310_7310.n493 w_13310_7310.n490 0.021
R606 w_13310_7310.n490 w_13310_7310.n488 0.021
R607 w_13310_7310.n488 w_13310_7310.n484 0.021
R608 w_13310_7310.n484 w_13310_7310.n482 0.021
R609 w_13310_7310.n482 w_13310_7310.n478 0.021
R610 w_13310_7310.n478 w_13310_7310.n476 0.021
R611 w_13310_7310.n476 w_13310_7310.n472 0.021
R612 w_13310_7310.n472 w_13310_7310.n470 0.021
R613 w_13310_7310.n470 w_13310_7310.n466 0.021
R614 w_13310_7310.n454 w_13310_7310.n452 0.021
R615 w_13310_7310.n452 w_13310_7310.n448 0.021
R616 w_13310_7310.n448 w_13310_7310.n446 0.021
R617 w_13310_7310.n446 w_13310_7310.n442 0.021
R618 w_13310_7310.n442 w_13310_7310.n440 0.021
R619 w_13310_7310.n440 w_13310_7310.n436 0.021
R620 w_13310_7310.n436 w_13310_7310.n434 0.021
R621 w_13310_7310.n434 w_13310_7310.n430 0.021
R622 w_13310_7310.n506 w_13310_7310.n503 0.021
R623 w_13310_7310.n508 w_13310_7310.n506 0.021
R624 w_13310_7310.n512 w_13310_7310.n508 0.021
R625 w_13310_7310.n514 w_13310_7310.n512 0.021
R626 w_13310_7310.n518 w_13310_7310.n514 0.021
R627 w_13310_7310.n520 w_13310_7310.n518 0.021
R628 w_13310_7310.n524 w_13310_7310.n520 0.021
R629 w_13310_7310.n526 w_13310_7310.n524 0.021
R630 w_13310_7310.n530 w_13310_7310.n526 0.021
R631 w_13310_7310.n532 w_13310_7310.n530 0.021
R632 w_13310_7310.n34 w_13310_7310.n32 0.021
R633 w_13310_7310.n32 w_13310_7310.n28 0.021
R634 w_13310_7310.n28 w_13310_7310.n26 0.021
R635 w_13310_7310.n26 w_13310_7310.n22 0.021
R636 w_13310_7310.n22 w_13310_7310.n20 0.021
R637 w_13310_7310.n20 w_13310_7310.n16 0.021
R638 w_13310_7310.n16 w_13310_7310.n14 0.021
R639 w_13310_7310.n14 w_13310_7310.n10 0.021
R640 w_13310_7310.n225 w_13310_7310.n221 0.021
R641 w_13310_7310.n301 w_13310_7310.n297 0.021
R642 w_13310_7310.n388 w_13310_7310.n384 0.021
R643 w_13310_7310.n464 w_13310_7310.n460 0.021
R644 w_13310_7310.n534 w_13310_7310.n533 0.021
R645 w_13310_7310.n146 w_13310_7310.n145 0.009
R646 w_13310_7310.n79 w_13310_7310.n78 0.009
R647 w_13310_7310.n221 w_13310_7310.n220 0.006
R648 w_13310_7310.n297 w_13310_7310.n296 0.006
R649 w_13310_7310.n384 w_13310_7310.n383 0.006
R650 w_13310_7310.n460 w_13310_7310.n459 0.006
R651 w_13310_7310.n534 w_13310_7310.n35 0.006
R652 a_800_7410.n7 a_800_7410.t22 708.072
R653 a_800_7410.n9 a_800_7410.t21 708.056
R654 a_800_7410.n11 a_800_7410.t14 708.054
R655 a_800_7410.n11 a_800_7410.t13 708.054
R656 a_800_7410.n9 a_800_7410.t17 708.05
R657 a_800_7410.n7 a_800_7410.t23 708.038
R658 a_800_7410.n6 a_800_7410.t16 388.574
R659 a_800_7410.n6 a_800_7410.t24 388.524
R660 a_800_7410.n12 a_800_7410.t18 388.509
R661 a_800_7410.n12 a_800_7410.t20 388.509
R662 a_800_7410.n10 a_800_7410.t19 388.509
R663 a_800_7410.n10 a_800_7410.t15 388.509
R664 a_800_7410.n13 a_800_7410.t0 5.713
R665 a_800_7410.n13 a_800_7410.t3 5.713
R666 a_800_7410.n5 a_800_7410.t6 5.713
R667 a_800_7410.n5 a_800_7410.t4 5.713
R668 a_800_7410.n3 a_800_7410.t2 5.713
R669 a_800_7410.n3 a_800_7410.t7 5.713
R670 a_800_7410.n4 a_800_7410.t8 3.48
R671 a_800_7410.n4 a_800_7410.t9 3.48
R672 a_800_7410.n2 a_800_7410.t5 3.48
R673 a_800_7410.n2 a_800_7410.t12 3.48
R674 a_800_7410.n14 a_800_7410.t11 3.48
R675 a_800_7410.t1 a_800_7410.n14 3.48
R676 a_800_7410.t10 a_800_7410.n1 2.751
R677 a_800_7410.n1 a_800_7410.n11 2.272
R678 a_800_7410.n8 a_800_7410.n7 2.265
R679 a_800_7410.n0 a_800_7410.n9 2.178
R680 a_800_7410.n5 a_800_7410.n4 1.164
R681 a_800_7410.n3 a_800_7410.n2 1.164
R682 a_800_7410.n14 a_800_7410.n13 1.112
R683 a_800_7410.n1 a_800_7410.n0 0.841
R684 a_800_7410.n0 a_800_7410.n8 0.804
R685 a_800_7410.n8 a_800_7410.n6 0.328
R686 a_800_7410.n1 a_800_7410.n12 0.29
R687 a_800_7410.t10 a_800_7410.n3 0.2
R688 a_800_7410.t10 a_800_7410.n5 0.2
R689 a_800_7410.n13 a_800_7410.t10 0.2
R690 a_800_7410.n0 a_800_7410.n10 0.162
R691 w_n4828_7260.n131 w_n4828_7260.t16 109.25
R692 w_n4828_7260.n173 w_n4828_7260.t14 109.25
R693 w_n4828_7260.n173 w_n4828_7260.t22 109.25
R694 w_n4828_7260.n225 w_n4828_7260.t10 109.25
R695 w_n4828_7260.n225 w_n4828_7260.t4 109.25
R696 w_n4828_7260.n288 w_n4828_7260.t34 109.25
R697 w_n4828_7260.n288 w_n4828_7260.t20 109.25
R698 w_n4828_7260.n362 w_n4828_7260.t2 109.25
R699 w_n4828_7260.n362 w_n4828_7260.t6 109.25
R700 w_n4828_7260.n396 w_n4828_7260.t32 109.25
R701 w_n4828_7260.n396 w_n4828_7260.t8 109.25
R702 w_n4828_7260.n94 w_n4828_7260.t0 109.25
R703 w_n4828_7260.n403 w_n4828_7260.n400 20.092
R704 w_n4828_7260.n99 w_n4828_7260.n98 16.607
R705 w_n4828_7260.n437 w_n4828_7260.n436 16.607
R706 w_n4828_7260.n339 w_n4828_7260.n338 16.289
R707 w_n4828_7260.n287 w_n4828_7260.n286 16.289
R708 w_n4828_7260.n224 w_n4828_7260.n223 16.289
R709 w_n4828_7260.n172 w_n4828_7260.n171 16.289
R710 w_n4828_7260.n75 w_n4828_7260.n71 12.923
R711 w_n4828_7260.n104 w_n4828_7260.n100 12.641
R712 w_n4828_7260.n181 w_n4828_7260.n177 12.629
R713 w_n4828_7260.n233 w_n4828_7260.n229 12.629
R714 w_n4828_7260.n296 w_n4828_7260.n292 12.629
R715 w_n4828_7260.n344 w_n4828_7260.n340 12.629
R716 w_n4828_7260.n106 w_n4828_7260.n105 9.3
R717 w_n4828_7260.n112 w_n4828_7260.n111 9.3
R718 w_n4828_7260.n118 w_n4828_7260.n117 9.3
R719 w_n4828_7260.n124 w_n4828_7260.n123 9.3
R720 w_n4828_7260.n130 w_n4828_7260.n129 9.3
R721 w_n4828_7260.n140 w_n4828_7260.n139 9.3
R722 w_n4828_7260.n146 w_n4828_7260.n145 9.3
R723 w_n4828_7260.n152 w_n4828_7260.n151 9.3
R724 w_n4828_7260.n158 w_n4828_7260.n157 9.3
R725 w_n4828_7260.n164 w_n4828_7260.n163 9.3
R726 w_n4828_7260.n169 w_n4828_7260.n168 9.3
R727 w_n4828_7260.n36 w_n4828_7260.n182 9.3
R728 w_n4828_7260.n35 w_n4828_7260.n186 9.3
R729 w_n4828_7260.n33 w_n4828_7260.n190 9.3
R730 w_n4828_7260.n34 w_n4828_7260.n194 9.3
R731 w_n4828_7260.n19 w_n4828_7260.n198 9.3
R732 w_n4828_7260.n0 w_n4828_7260.n202 9.3
R733 w_n4828_7260.n32 w_n4828_7260.n206 9.3
R734 w_n4828_7260.n31 w_n4828_7260.n210 9.3
R735 w_n4828_7260.n30 w_n4828_7260.n214 9.3
R736 w_n4828_7260.n20 w_n4828_7260.n218 9.3
R737 w_n4828_7260.n21 w_n4828_7260.n221 9.3
R738 w_n4828_7260.n43 w_n4828_7260.n234 9.3
R739 w_n4828_7260.n42 w_n4828_7260.n238 9.3
R740 w_n4828_7260.n40 w_n4828_7260.n242 9.3
R741 w_n4828_7260.n41 w_n4828_7260.n246 9.3
R742 w_n4828_7260.n18 w_n4828_7260.n250 9.3
R743 w_n4828_7260.n1 w_n4828_7260.n254 9.3
R744 w_n4828_7260.n39 w_n4828_7260.n258 9.3
R745 w_n4828_7260.n38 w_n4828_7260.n262 9.3
R746 w_n4828_7260.n37 w_n4828_7260.n266 9.3
R747 w_n4828_7260.n22 w_n4828_7260.n270 9.3
R748 w_n4828_7260.n23 w_n4828_7260.n273 9.3
R749 w_n4828_7260.n50 w_n4828_7260.n297 9.3
R750 w_n4828_7260.n49 w_n4828_7260.n301 9.3
R751 w_n4828_7260.n47 w_n4828_7260.n305 9.3
R752 w_n4828_7260.n48 w_n4828_7260.n309 9.3
R753 w_n4828_7260.n17 w_n4828_7260.n313 9.3
R754 w_n4828_7260.n2 w_n4828_7260.n317 9.3
R755 w_n4828_7260.n46 w_n4828_7260.n321 9.3
R756 w_n4828_7260.n45 w_n4828_7260.n325 9.3
R757 w_n4828_7260.n44 w_n4828_7260.n329 9.3
R758 w_n4828_7260.n24 w_n4828_7260.n333 9.3
R759 w_n4828_7260.n25 w_n4828_7260.n336 9.3
R760 w_n4828_7260.n57 w_n4828_7260.n345 9.3
R761 w_n4828_7260.n56 w_n4828_7260.n349 9.3
R762 w_n4828_7260.n54 w_n4828_7260.n353 9.3
R763 w_n4828_7260.n55 w_n4828_7260.n357 9.3
R764 w_n4828_7260.n16 w_n4828_7260.n361 9.3
R765 w_n4828_7260.n3 w_n4828_7260.n369 9.3
R766 w_n4828_7260.n53 w_n4828_7260.n373 9.3
R767 w_n4828_7260.n52 w_n4828_7260.n377 9.3
R768 w_n4828_7260.n51 w_n4828_7260.n381 9.3
R769 w_n4828_7260.n26 w_n4828_7260.n385 9.3
R770 w_n4828_7260.n27 w_n4828_7260.n388 9.3
R771 w_n4828_7260.n57 w_n4828_7260.n348 9.3
R772 w_n4828_7260.n56 w_n4828_7260.n352 9.3
R773 w_n4828_7260.n54 w_n4828_7260.n356 9.3
R774 w_n4828_7260.n55 w_n4828_7260.n360 9.3
R775 w_n4828_7260.n3 w_n4828_7260.n372 9.3
R776 w_n4828_7260.n53 w_n4828_7260.n376 9.3
R777 w_n4828_7260.n52 w_n4828_7260.n380 9.3
R778 w_n4828_7260.n51 w_n4828_7260.n384 9.3
R779 w_n4828_7260.n26 w_n4828_7260.n387 9.3
R780 w_n4828_7260.n50 w_n4828_7260.n300 9.3
R781 w_n4828_7260.n49 w_n4828_7260.n304 9.3
R782 w_n4828_7260.n47 w_n4828_7260.n308 9.3
R783 w_n4828_7260.n48 w_n4828_7260.n312 9.3
R784 w_n4828_7260.n2 w_n4828_7260.n320 9.3
R785 w_n4828_7260.n46 w_n4828_7260.n324 9.3
R786 w_n4828_7260.n45 w_n4828_7260.n328 9.3
R787 w_n4828_7260.n44 w_n4828_7260.n332 9.3
R788 w_n4828_7260.n24 w_n4828_7260.n335 9.3
R789 w_n4828_7260.n43 w_n4828_7260.n237 9.3
R790 w_n4828_7260.n42 w_n4828_7260.n241 9.3
R791 w_n4828_7260.n40 w_n4828_7260.n245 9.3
R792 w_n4828_7260.n41 w_n4828_7260.n249 9.3
R793 w_n4828_7260.n1 w_n4828_7260.n257 9.3
R794 w_n4828_7260.n39 w_n4828_7260.n261 9.3
R795 w_n4828_7260.n38 w_n4828_7260.n265 9.3
R796 w_n4828_7260.n37 w_n4828_7260.n269 9.3
R797 w_n4828_7260.n22 w_n4828_7260.n272 9.3
R798 w_n4828_7260.n36 w_n4828_7260.n185 9.3
R799 w_n4828_7260.n35 w_n4828_7260.n189 9.3
R800 w_n4828_7260.n33 w_n4828_7260.n193 9.3
R801 w_n4828_7260.n34 w_n4828_7260.n197 9.3
R802 w_n4828_7260.n0 w_n4828_7260.n205 9.3
R803 w_n4828_7260.n32 w_n4828_7260.n209 9.3
R804 w_n4828_7260.n31 w_n4828_7260.n213 9.3
R805 w_n4828_7260.n30 w_n4828_7260.n217 9.3
R806 w_n4828_7260.n20 w_n4828_7260.n220 9.3
R807 w_n4828_7260.n110 w_n4828_7260.n109 9.3
R808 w_n4828_7260.n116 w_n4828_7260.n115 9.3
R809 w_n4828_7260.n122 w_n4828_7260.n121 9.3
R810 w_n4828_7260.n128 w_n4828_7260.n127 9.3
R811 w_n4828_7260.n144 w_n4828_7260.n143 9.3
R812 w_n4828_7260.n150 w_n4828_7260.n149 9.3
R813 w_n4828_7260.n156 w_n4828_7260.n155 9.3
R814 w_n4828_7260.n162 w_n4828_7260.n161 9.3
R815 w_n4828_7260.n167 w_n4828_7260.n166 9.3
R816 w_n4828_7260.n64 w_n4828_7260.n404 9.3
R817 w_n4828_7260.n64 w_n4828_7260.n406 9.3
R818 w_n4828_7260.n63 w_n4828_7260.n407 9.3
R819 w_n4828_7260.n63 w_n4828_7260.n409 9.3
R820 w_n4828_7260.n61 w_n4828_7260.n410 9.3
R821 w_n4828_7260.n61 w_n4828_7260.n412 9.3
R822 w_n4828_7260.n62 w_n4828_7260.n413 9.3
R823 w_n4828_7260.n62 w_n4828_7260.n415 9.3
R824 w_n4828_7260.n15 w_n4828_7260.n416 9.3
R825 w_n4828_7260.n4 w_n4828_7260.n419 9.3
R826 w_n4828_7260.n4 w_n4828_7260.n421 9.3
R827 w_n4828_7260.n60 w_n4828_7260.n422 9.3
R828 w_n4828_7260.n60 w_n4828_7260.n424 9.3
R829 w_n4828_7260.n59 w_n4828_7260.n425 9.3
R830 w_n4828_7260.n59 w_n4828_7260.n427 9.3
R831 w_n4828_7260.n58 w_n4828_7260.n428 9.3
R832 w_n4828_7260.n58 w_n4828_7260.n430 9.3
R833 w_n4828_7260.n28 w_n4828_7260.n431 9.3
R834 w_n4828_7260.n28 w_n4828_7260.n433 9.3
R835 w_n4828_7260.n29 w_n4828_7260.n434 9.3
R836 w_n4828_7260.n5 w_n4828_7260.n439 9.3
R837 w_n4828_7260.n14 w_n4828_7260.n76 9.3
R838 w_n4828_7260.n14 w_n4828_7260.n79 9.3
R839 w_n4828_7260.n13 w_n4828_7260.n80 9.3
R840 w_n4828_7260.n13 w_n4828_7260.n83 9.3
R841 w_n4828_7260.n11 w_n4828_7260.n84 9.3
R842 w_n4828_7260.n11 w_n4828_7260.n87 9.3
R843 w_n4828_7260.n12 w_n4828_7260.n88 9.3
R844 w_n4828_7260.n12 w_n4828_7260.n91 9.3
R845 w_n4828_7260.n93 w_n4828_7260.n92 9.3
R846 w_n4828_7260.n10 w_n4828_7260.n458 9.3
R847 w_n4828_7260.n10 w_n4828_7260.n457 9.3
R848 w_n4828_7260.n9 w_n4828_7260.n454 9.3
R849 w_n4828_7260.n9 w_n4828_7260.n453 9.3
R850 w_n4828_7260.n8 w_n4828_7260.n450 9.3
R851 w_n4828_7260.n8 w_n4828_7260.n449 9.3
R852 w_n4828_7260.n7 w_n4828_7260.n446 9.3
R853 w_n4828_7260.n7 w_n4828_7260.n445 9.3
R854 w_n4828_7260.n6 w_n4828_7260.n442 9.3
R855 w_n4828_7260.n6 w_n4828_7260.n441 9.3
R856 w_n4828_7260.n343 w_n4828_7260.n342 8.855
R857 w_n4828_7260.n348 w_n4828_7260.n347 8.855
R858 w_n4828_7260.n352 w_n4828_7260.n351 8.855
R859 w_n4828_7260.n356 w_n4828_7260.n355 8.855
R860 w_n4828_7260.n360 w_n4828_7260.n359 8.855
R861 w_n4828_7260.n365 w_n4828_7260.n364 8.855
R862 w_n4828_7260.n368 w_n4828_7260.n367 8.855
R863 w_n4828_7260.n372 w_n4828_7260.n371 8.855
R864 w_n4828_7260.n376 w_n4828_7260.n375 8.855
R865 w_n4828_7260.n380 w_n4828_7260.n379 8.855
R866 w_n4828_7260.n384 w_n4828_7260.n383 8.855
R867 w_n4828_7260.n387 w_n4828_7260.n386 8.855
R868 w_n4828_7260.n295 w_n4828_7260.n294 8.855
R869 w_n4828_7260.n300 w_n4828_7260.n299 8.855
R870 w_n4828_7260.n304 w_n4828_7260.n303 8.855
R871 w_n4828_7260.n308 w_n4828_7260.n307 8.855
R872 w_n4828_7260.n312 w_n4828_7260.n311 8.855
R873 w_n4828_7260.n291 w_n4828_7260.n290 8.855
R874 w_n4828_7260.n316 w_n4828_7260.n315 8.855
R875 w_n4828_7260.n320 w_n4828_7260.n319 8.855
R876 w_n4828_7260.n324 w_n4828_7260.n323 8.855
R877 w_n4828_7260.n328 w_n4828_7260.n327 8.855
R878 w_n4828_7260.n332 w_n4828_7260.n331 8.855
R879 w_n4828_7260.n335 w_n4828_7260.n334 8.855
R880 w_n4828_7260.n232 w_n4828_7260.n231 8.855
R881 w_n4828_7260.n237 w_n4828_7260.n236 8.855
R882 w_n4828_7260.n241 w_n4828_7260.n240 8.855
R883 w_n4828_7260.n245 w_n4828_7260.n244 8.855
R884 w_n4828_7260.n249 w_n4828_7260.n248 8.855
R885 w_n4828_7260.n228 w_n4828_7260.n227 8.855
R886 w_n4828_7260.n253 w_n4828_7260.n252 8.855
R887 w_n4828_7260.n257 w_n4828_7260.n256 8.855
R888 w_n4828_7260.n261 w_n4828_7260.n260 8.855
R889 w_n4828_7260.n265 w_n4828_7260.n264 8.855
R890 w_n4828_7260.n269 w_n4828_7260.n268 8.855
R891 w_n4828_7260.n272 w_n4828_7260.n271 8.855
R892 w_n4828_7260.n180 w_n4828_7260.n179 8.855
R893 w_n4828_7260.n185 w_n4828_7260.n184 8.855
R894 w_n4828_7260.n189 w_n4828_7260.n188 8.855
R895 w_n4828_7260.n193 w_n4828_7260.n192 8.855
R896 w_n4828_7260.n197 w_n4828_7260.n196 8.855
R897 w_n4828_7260.n176 w_n4828_7260.n175 8.855
R898 w_n4828_7260.n201 w_n4828_7260.n200 8.855
R899 w_n4828_7260.n205 w_n4828_7260.n204 8.855
R900 w_n4828_7260.n209 w_n4828_7260.n208 8.855
R901 w_n4828_7260.n213 w_n4828_7260.n212 8.855
R902 w_n4828_7260.n217 w_n4828_7260.n216 8.855
R903 w_n4828_7260.n220 w_n4828_7260.n219 8.855
R904 w_n4828_7260.n103 w_n4828_7260.n102 8.855
R905 w_n4828_7260.n109 w_n4828_7260.n108 8.855
R906 w_n4828_7260.n115 w_n4828_7260.n114 8.855
R907 w_n4828_7260.n121 w_n4828_7260.n120 8.855
R908 w_n4828_7260.n127 w_n4828_7260.n126 8.855
R909 w_n4828_7260.n134 w_n4828_7260.n133 8.855
R910 w_n4828_7260.n137 w_n4828_7260.n136 8.855
R911 w_n4828_7260.n143 w_n4828_7260.n142 8.855
R912 w_n4828_7260.n149 w_n4828_7260.n148 8.855
R913 w_n4828_7260.n155 w_n4828_7260.n154 8.855
R914 w_n4828_7260.n161 w_n4828_7260.n160 8.855
R915 w_n4828_7260.n166 w_n4828_7260.n165 8.855
R916 w_n4828_7260.n74 w_n4828_7260.n73 8.855
R917 w_n4828_7260.n402 w_n4828_7260.n401 8.855
R918 w_n4828_7260.n406 w_n4828_7260.n405 8.855
R919 w_n4828_7260.n409 w_n4828_7260.n408 8.855
R920 w_n4828_7260.n412 w_n4828_7260.n411 8.855
R921 w_n4828_7260.n415 w_n4828_7260.n414 8.855
R922 w_n4828_7260.n399 w_n4828_7260.n398 8.855
R923 w_n4828_7260.n418 w_n4828_7260.n417 8.855
R924 w_n4828_7260.n421 w_n4828_7260.n420 8.855
R925 w_n4828_7260.n424 w_n4828_7260.n423 8.855
R926 w_n4828_7260.n427 w_n4828_7260.n426 8.855
R927 w_n4828_7260.n430 w_n4828_7260.n429 8.855
R928 w_n4828_7260.n433 w_n4828_7260.n432 8.855
R929 w_n4828_7260.n79 w_n4828_7260.n78 8.855
R930 w_n4828_7260.n83 w_n4828_7260.n82 8.855
R931 w_n4828_7260.n87 w_n4828_7260.n86 8.855
R932 w_n4828_7260.n91 w_n4828_7260.n90 8.855
R933 w_n4828_7260.n70 w_n4828_7260.n69 8.855
R934 w_n4828_7260.n97 w_n4828_7260.n96 8.855
R935 w_n4828_7260.n457 w_n4828_7260.n456 8.855
R936 w_n4828_7260.n453 w_n4828_7260.n452 8.855
R937 w_n4828_7260.n449 w_n4828_7260.n448 8.855
R938 w_n4828_7260.n445 w_n4828_7260.n444 8.855
R939 w_n4828_7260.n441 w_n4828_7260.n440 8.855
R940 w_n4828_7260.n398 w_n4828_7260.n397 7.463
R941 w_n4828_7260.n27 w_n4828_7260.n339 6.209
R942 w_n4828_7260.n25 w_n4828_7260.n287 6.209
R943 w_n4828_7260.n23 w_n4828_7260.n224 6.209
R944 w_n4828_7260.n21 w_n4828_7260.n172 6.209
R945 w_n4828_7260.n29 w_n4828_7260.n390 6.209
R946 w_n4828_7260.n170 w_n4828_7260.n99 6.208
R947 w_n4828_7260.n363 w_n4828_7260.n362 5.95
R948 w_n4828_7260.n289 w_n4828_7260.n288 5.95
R949 w_n4828_7260.n226 w_n4828_7260.n225 5.95
R950 w_n4828_7260.n174 w_n4828_7260.n173 5.95
R951 w_n4828_7260.n3 w_n4828_7260.n368 5.876
R952 w_n4828_7260.n2 w_n4828_7260.n316 5.876
R953 w_n4828_7260.n1 w_n4828_7260.n253 5.876
R954 w_n4828_7260.n0 w_n4828_7260.n201 5.876
R955 w_n4828_7260.n4 w_n4828_7260.n418 5.876
R956 w_n4828_7260.n65 w_n4828_7260.n70 5.873
R957 w_n4828_7260.n138 w_n4828_7260.n137 5.873
R958 w_n4828_7260.n4 w_n4828_7260.t33 5.713
R959 w_n4828_7260.n3 w_n4828_7260.t3 5.713
R960 w_n4828_7260.n3 w_n4828_7260.t7 5.713
R961 w_n4828_7260.n67 w_n4828_7260.t17 5.713
R962 w_n4828_7260.n0 w_n4828_7260.t15 5.713
R963 w_n4828_7260.n0 w_n4828_7260.t23 5.713
R964 w_n4828_7260.n1 w_n4828_7260.t11 5.713
R965 w_n4828_7260.n1 w_n4828_7260.t5 5.713
R966 w_n4828_7260.n2 w_n4828_7260.t35 5.713
R967 w_n4828_7260.n2 w_n4828_7260.t21 5.713
R968 w_n4828_7260.n4 w_n4828_7260.t9 5.713
R969 w_n4828_7260.t1 w_n4828_7260.n66 5.713
R970 w_n4828_7260.n438 w_n4828_7260.n437 5.637
R971 w_n4828_7260.n181 w_n4828_7260.n180 5.614
R972 w_n4828_7260.n233 w_n4828_7260.n232 5.614
R973 w_n4828_7260.n296 w_n4828_7260.n295 5.614
R974 w_n4828_7260.n344 w_n4828_7260.n343 5.614
R975 w_n4828_7260.n403 w_n4828_7260.n402 5.614
R976 w_n4828_7260.n104 w_n4828_7260.n103 5.611
R977 w_n4828_7260.n75 w_n4828_7260.n74 5.571
R978 w_n4828_7260.n132 w_n4828_7260.n131 5.347
R979 w_n4828_7260.n95 w_n4828_7260.n94 5.347
R980 w_n4828_7260.n275 w_n4828_7260.t27 4.491
R981 w_n4828_7260.n275 w_n4828_7260.t29 4.386
R982 w_n4828_7260.n276 w_n4828_7260.t18 4.386
R983 w_n4828_7260.n277 w_n4828_7260.t19 4.386
R984 w_n4828_7260.n278 w_n4828_7260.t28 4.386
R985 w_n4828_7260.n279 w_n4828_7260.t31 4.386
R986 w_n4828_7260.n280 w_n4828_7260.t13 4.386
R987 w_n4828_7260.n281 w_n4828_7260.t25 4.386
R988 w_n4828_7260.n282 w_n4828_7260.t30 4.386
R989 w_n4828_7260.n283 w_n4828_7260.t26 4.386
R990 w_n4828_7260.n284 w_n4828_7260.t24 4.386
R991 w_n4828_7260.n285 w_n4828_7260.t12 4.386
R992 w_n4828_7260.n3 w_n4828_7260.n365 4.27
R993 w_n4828_7260.n2 w_n4828_7260.n291 4.27
R994 w_n4828_7260.n1 w_n4828_7260.n228 4.27
R995 w_n4828_7260.n0 w_n4828_7260.n176 4.27
R996 w_n4828_7260.n4 w_n4828_7260.n399 4.27
R997 w_n4828_7260.n67 w_n4828_7260.n134 4.269
R998 w_n4828_7260.n66 w_n4828_7260.n97 4.269
R999 w_n4828_7260.n444 w_n4828_7260.n443 3.685
R1000 w_n4828_7260.n448 w_n4828_7260.n447 3.685
R1001 w_n4828_7260.n452 w_n4828_7260.n451 3.685
R1002 w_n4828_7260.n456 w_n4828_7260.n455 3.685
R1003 w_n4828_7260.n96 w_n4828_7260.n95 3.685
R1004 w_n4828_7260.n69 w_n4828_7260.n68 3.685
R1005 w_n4828_7260.n90 w_n4828_7260.n89 3.685
R1006 w_n4828_7260.n86 w_n4828_7260.n85 3.685
R1007 w_n4828_7260.n82 w_n4828_7260.n81 3.685
R1008 w_n4828_7260.n78 w_n4828_7260.n77 3.685
R1009 w_n4828_7260.n160 w_n4828_7260.n159 3.685
R1010 w_n4828_7260.n154 w_n4828_7260.n153 3.685
R1011 w_n4828_7260.n148 w_n4828_7260.n147 3.685
R1012 w_n4828_7260.n142 w_n4828_7260.n141 3.685
R1013 w_n4828_7260.n136 w_n4828_7260.n135 3.685
R1014 w_n4828_7260.n133 w_n4828_7260.n132 3.685
R1015 w_n4828_7260.n126 w_n4828_7260.n125 3.685
R1016 w_n4828_7260.n120 w_n4828_7260.n119 3.685
R1017 w_n4828_7260.n114 w_n4828_7260.n113 3.685
R1018 w_n4828_7260.n108 w_n4828_7260.n107 3.685
R1019 w_n4828_7260.n73 w_n4828_7260.n72 3.514
R1020 w_n4828_7260.n102 w_n4828_7260.n101 3.514
R1021 w_n4828_7260.n216 w_n4828_7260.n215 3.052
R1022 w_n4828_7260.n212 w_n4828_7260.n211 3.052
R1023 w_n4828_7260.n208 w_n4828_7260.n207 3.052
R1024 w_n4828_7260.n204 w_n4828_7260.n203 3.052
R1025 w_n4828_7260.n200 w_n4828_7260.n199 3.052
R1026 w_n4828_7260.n175 w_n4828_7260.n174 3.052
R1027 w_n4828_7260.n196 w_n4828_7260.n195 3.052
R1028 w_n4828_7260.n192 w_n4828_7260.n191 3.052
R1029 w_n4828_7260.n188 w_n4828_7260.n187 3.052
R1030 w_n4828_7260.n184 w_n4828_7260.n183 3.052
R1031 w_n4828_7260.n268 w_n4828_7260.n267 3.052
R1032 w_n4828_7260.n264 w_n4828_7260.n263 3.052
R1033 w_n4828_7260.n260 w_n4828_7260.n259 3.052
R1034 w_n4828_7260.n256 w_n4828_7260.n255 3.052
R1035 w_n4828_7260.n252 w_n4828_7260.n251 3.052
R1036 w_n4828_7260.n227 w_n4828_7260.n226 3.052
R1037 w_n4828_7260.n248 w_n4828_7260.n247 3.052
R1038 w_n4828_7260.n244 w_n4828_7260.n243 3.052
R1039 w_n4828_7260.n240 w_n4828_7260.n239 3.052
R1040 w_n4828_7260.n236 w_n4828_7260.n235 3.052
R1041 w_n4828_7260.n331 w_n4828_7260.n330 3.052
R1042 w_n4828_7260.n327 w_n4828_7260.n326 3.052
R1043 w_n4828_7260.n323 w_n4828_7260.n322 3.052
R1044 w_n4828_7260.n319 w_n4828_7260.n318 3.052
R1045 w_n4828_7260.n315 w_n4828_7260.n314 3.052
R1046 w_n4828_7260.n290 w_n4828_7260.n289 3.052
R1047 w_n4828_7260.n311 w_n4828_7260.n310 3.052
R1048 w_n4828_7260.n307 w_n4828_7260.n306 3.052
R1049 w_n4828_7260.n303 w_n4828_7260.n302 3.052
R1050 w_n4828_7260.n299 w_n4828_7260.n298 3.052
R1051 w_n4828_7260.n383 w_n4828_7260.n382 3.052
R1052 w_n4828_7260.n379 w_n4828_7260.n378 3.052
R1053 w_n4828_7260.n375 w_n4828_7260.n374 3.052
R1054 w_n4828_7260.n371 w_n4828_7260.n370 3.052
R1055 w_n4828_7260.n367 w_n4828_7260.n366 3.052
R1056 w_n4828_7260.n364 w_n4828_7260.n363 3.052
R1057 w_n4828_7260.n359 w_n4828_7260.n358 3.052
R1058 w_n4828_7260.n355 w_n4828_7260.n354 3.052
R1059 w_n4828_7260.n351 w_n4828_7260.n350 3.052
R1060 w_n4828_7260.n347 w_n4828_7260.n346 3.052
R1061 w_n4828_7260.n179 w_n4828_7260.n178 2.91
R1062 w_n4828_7260.n231 w_n4828_7260.n230 2.91
R1063 w_n4828_7260.n294 w_n4828_7260.n293 2.91
R1064 w_n4828_7260.n342 w_n4828_7260.n341 2.91
R1065 w_n4828_7260.n337 w_n4828_7260.n285 2.206
R1066 w_n4828_7260.n438 w_n4828_7260.n435 0.768
R1067 w_n4828_7260.n222 w_n4828_7260.n170 0.75
R1068 w_n4828_7260.n14 w_n4828_7260.n75 0.713
R1069 w_n4828_7260.n396 w_n4828_7260.n395 0.697
R1070 w_n4828_7260.n396 w_n4828_7260.n394 0.697
R1071 w_n4828_7260.n397 w_n4828_7260.n396 0.697
R1072 w_n4828_7260.n396 w_n4828_7260.n393 0.697
R1073 w_n4828_7260.n396 w_n4828_7260.n392 0.697
R1074 w_n4828_7260.n396 w_n4828_7260.n391 0.697
R1075 w_n4828_7260.n106 w_n4828_7260.n104 0.668
R1076 w_n4828_7260.n64 w_n4828_7260.n403 0.652
R1077 w_n4828_7260.n36 w_n4828_7260.n181 0.652
R1078 w_n4828_7260.n43 w_n4828_7260.n233 0.652
R1079 w_n4828_7260.n50 w_n4828_7260.n296 0.652
R1080 w_n4828_7260.n57 w_n4828_7260.n344 0.652
R1081 w_n4828_7260.n274 w_n4828_7260.n222 0.57
R1082 w_n4828_7260.n337 w_n4828_7260.n274 0.57
R1083 w_n4828_7260.n435 w_n4828_7260.n389 0.57
R1084 w_n4828_7260.n389 w_n4828_7260.n337 0.57
R1085 w_n4828_7260.n222 w_n4828_7260.n21 0.208
R1086 w_n4828_7260.n274 w_n4828_7260.n23 0.208
R1087 w_n4828_7260.n337 w_n4828_7260.n25 0.208
R1088 w_n4828_7260.n389 w_n4828_7260.n27 0.208
R1089 w_n4828_7260.n435 w_n4828_7260.n29 0.208
R1090 w_n4828_7260.n277 w_n4828_7260.n276 0.106
R1091 w_n4828_7260.n279 w_n4828_7260.n278 0.106
R1092 w_n4828_7260.n281 w_n4828_7260.n280 0.106
R1093 w_n4828_7260.n283 w_n4828_7260.n282 0.106
R1094 w_n4828_7260.n285 w_n4828_7260.n284 0.106
R1095 w_n4828_7260.n276 w_n4828_7260.n275 0.083
R1096 w_n4828_7260.n278 w_n4828_7260.n277 0.083
R1097 w_n4828_7260.n280 w_n4828_7260.n279 0.083
R1098 w_n4828_7260.n282 w_n4828_7260.n281 0.083
R1099 w_n4828_7260.n284 w_n4828_7260.n283 0.083
R1100 w_n4828_7260.n60 w_n4828_7260.n4 0.073
R1101 w_n4828_7260.n53 w_n4828_7260.n3 0.073
R1102 w_n4828_7260.n46 w_n4828_7260.n2 0.073
R1103 w_n4828_7260.n39 w_n4828_7260.n1 0.073
R1104 w_n4828_7260.n32 w_n4828_7260.n0 0.073
R1105 w_n4828_7260.n29 w_n4828_7260.n28 0.069
R1106 w_n4828_7260.n27 w_n4828_7260.n26 0.069
R1107 w_n4828_7260.n25 w_n4828_7260.n24 0.069
R1108 w_n4828_7260.n23 w_n4828_7260.n22 0.069
R1109 w_n4828_7260.n21 w_n4828_7260.n20 0.069
R1110 w_n4828_7260.n13 w_n4828_7260.n14 0.062
R1111 w_n4828_7260.n11 w_n4828_7260.n13 0.062
R1112 w_n4828_7260.n12 w_n4828_7260.n11 0.062
R1113 w_n4828_7260.n93 w_n4828_7260.n12 0.062
R1114 w_n4828_7260.n10 w_n4828_7260.n9 0.062
R1115 w_n4828_7260.n9 w_n4828_7260.n8 0.062
R1116 w_n4828_7260.n8 w_n4828_7260.n7 0.062
R1117 w_n4828_7260.n7 w_n4828_7260.n6 0.062
R1118 w_n4828_7260.n6 w_n4828_7260.n5 0.062
R1119 w_n4828_7260.n0 w_n4828_7260.n19 0.056
R1120 w_n4828_7260.n1 w_n4828_7260.n18 0.056
R1121 w_n4828_7260.n2 w_n4828_7260.n17 0.056
R1122 w_n4828_7260.n3 w_n4828_7260.n16 0.056
R1123 w_n4828_7260.n4 w_n4828_7260.n15 0.056
R1124 w_n4828_7260.n140 w_n4828_7260.n138 0.047
R1125 w_n4828_7260.n65 w_n4828_7260.n93 0.046
R1126 w_n4828_7260.n5 w_n4828_7260.n438 0.045
R1127 w_n4828_7260.n67 w_n4828_7260.n130 0.043
R1128 w_n4828_7260.n63 w_n4828_7260.n64 0.042
R1129 w_n4828_7260.n61 w_n4828_7260.n63 0.042
R1130 w_n4828_7260.n62 w_n4828_7260.n61 0.042
R1131 w_n4828_7260.n15 w_n4828_7260.n62 0.042
R1132 w_n4828_7260.n59 w_n4828_7260.n60 0.042
R1133 w_n4828_7260.n58 w_n4828_7260.n59 0.042
R1134 w_n4828_7260.n28 w_n4828_7260.n58 0.042
R1135 w_n4828_7260.n56 w_n4828_7260.n57 0.042
R1136 w_n4828_7260.n54 w_n4828_7260.n56 0.042
R1137 w_n4828_7260.n55 w_n4828_7260.n54 0.042
R1138 w_n4828_7260.n16 w_n4828_7260.n55 0.042
R1139 w_n4828_7260.n52 w_n4828_7260.n53 0.042
R1140 w_n4828_7260.n51 w_n4828_7260.n52 0.042
R1141 w_n4828_7260.n26 w_n4828_7260.n51 0.042
R1142 w_n4828_7260.n49 w_n4828_7260.n50 0.042
R1143 w_n4828_7260.n47 w_n4828_7260.n49 0.042
R1144 w_n4828_7260.n48 w_n4828_7260.n47 0.042
R1145 w_n4828_7260.n17 w_n4828_7260.n48 0.042
R1146 w_n4828_7260.n45 w_n4828_7260.n46 0.042
R1147 w_n4828_7260.n44 w_n4828_7260.n45 0.042
R1148 w_n4828_7260.n24 w_n4828_7260.n44 0.042
R1149 w_n4828_7260.n42 w_n4828_7260.n43 0.042
R1150 w_n4828_7260.n40 w_n4828_7260.n42 0.042
R1151 w_n4828_7260.n41 w_n4828_7260.n40 0.042
R1152 w_n4828_7260.n18 w_n4828_7260.n41 0.042
R1153 w_n4828_7260.n38 w_n4828_7260.n39 0.042
R1154 w_n4828_7260.n37 w_n4828_7260.n38 0.042
R1155 w_n4828_7260.n22 w_n4828_7260.n37 0.042
R1156 w_n4828_7260.n35 w_n4828_7260.n36 0.042
R1157 w_n4828_7260.n33 w_n4828_7260.n35 0.042
R1158 w_n4828_7260.n34 w_n4828_7260.n33 0.042
R1159 w_n4828_7260.n19 w_n4828_7260.n34 0.042
R1160 w_n4828_7260.n31 w_n4828_7260.n32 0.042
R1161 w_n4828_7260.n30 w_n4828_7260.n31 0.042
R1162 w_n4828_7260.n20 w_n4828_7260.n30 0.042
R1163 w_n4828_7260.n66 w_n4828_7260.n10 0.042
R1164 w_n4828_7260.n170 w_n4828_7260.n169 0.04
R1165 w_n4828_7260.n138 w_n4828_7260.n67 0.04
R1166 w_n4828_7260.n66 w_n4828_7260.n65 0.039
R1167 w_n4828_7260.n169 w_n4828_7260.n167 0.032
R1168 w_n4828_7260.n167 w_n4828_7260.n164 0.032
R1169 w_n4828_7260.n164 w_n4828_7260.n162 0.032
R1170 w_n4828_7260.n162 w_n4828_7260.n158 0.032
R1171 w_n4828_7260.n158 w_n4828_7260.n156 0.032
R1172 w_n4828_7260.n156 w_n4828_7260.n152 0.032
R1173 w_n4828_7260.n152 w_n4828_7260.n150 0.032
R1174 w_n4828_7260.n150 w_n4828_7260.n146 0.032
R1175 w_n4828_7260.n146 w_n4828_7260.n144 0.032
R1176 w_n4828_7260.n144 w_n4828_7260.n140 0.032
R1177 w_n4828_7260.n130 w_n4828_7260.n128 0.032
R1178 w_n4828_7260.n128 w_n4828_7260.n124 0.032
R1179 w_n4828_7260.n124 w_n4828_7260.n122 0.032
R1180 w_n4828_7260.n122 w_n4828_7260.n118 0.032
R1181 w_n4828_7260.n118 w_n4828_7260.n116 0.032
R1182 w_n4828_7260.n116 w_n4828_7260.n112 0.032
R1183 w_n4828_7260.n112 w_n4828_7260.n110 0.032
R1184 w_n4828_7260.n110 w_n4828_7260.n106 0.032
R1185 a_730_7313.n8 a_730_7313.t19 708.034
R1186 a_730_7313.n7 a_730_7313.t21 708.034
R1187 a_730_7313.n10 a_730_7313.t23 708.034
R1188 a_730_7313.n8 a_730_7313.t22 708.034
R1189 a_730_7313.n7 a_730_7313.t15 708.034
R1190 a_730_7313.n10 a_730_7313.t24 708.034
R1191 a_730_7313.n11 a_730_7313.t14 388.664
R1192 a_730_7313.n9 a_730_7313.t18 388.587
R1193 a_730_7313.n9 a_730_7313.t13 388.587
R1194 a_730_7313.n6 a_730_7313.t12 388.587
R1195 a_730_7313.n6 a_730_7313.t20 388.587
R1196 a_730_7313.n11 a_730_7313.t16 388.543
R1197 a_730_7313.n18 a_730_7313.t11 5.713
R1198 a_730_7313.n18 a_730_7313.t8 5.713
R1199 a_730_7313.n3 a_730_7313.t7 5.713
R1200 a_730_7313.n3 a_730_7313.t10 5.713
R1201 a_730_7313.n15 a_730_7313.t0 5.713
R1202 a_730_7313.n15 a_730_7313.t9 5.713
R1203 a_730_7313.n2 a_730_7313.t1 3.48
R1204 a_730_7313.n2 a_730_7313.t2 3.48
R1205 a_730_7313.n14 a_730_7313.t4 3.48
R1206 a_730_7313.n14 a_730_7313.t3 3.48
R1207 a_730_7313.n20 a_730_7313.t5 3.48
R1208 a_730_7313.t6 a_730_7313.n20 3.48
R1209 a_730_7313.n13 a_730_7313.n0 2.556
R1210 a_730_7313.n0 a_730_7313.n7 2.489
R1211 a_730_7313.n12 a_730_7313.n10 2.478
R1212 a_730_7313.n1 a_730_7313.n8 2.348
R1213 a_730_7313.n0 a_730_7313.n1 0.841
R1214 a_730_7313.n1 a_730_7313.n12 0.819
R1215 a_730_7313.n4 a_730_7313.n2 0.701
R1216 a_730_7313.n16 a_730_7313.n14 0.701
R1217 a_730_7313.n20 a_730_7313.n19 0.701
R1218 a_730_7313.n16 a_730_7313.n15 0.463
R1219 a_730_7313.n19 a_730_7313.n18 0.463
R1220 a_730_7313.n4 a_730_7313.n3 0.419
R1221 a_730_7313.n19 a_730_7313.t17 0.141
R1222 a_730_7313.n17 a_730_7313.n16 0.116
R1223 a_730_7313.t17 a_730_7313.n17 0.115
R1224 a_730_7313.n5 a_730_7313.n4 0.112
R1225 a_730_7313.n12 a_730_7313.n11 0.099
R1226 a_730_7313.n0 a_730_7313.n6 0.077
R1227 a_730_7313.n13 a_730_7313.n5 0.058
R1228 a_730_7313.n1 a_730_7313.n9 0.03
R1229 a_730_7313.t17 a_730_7313.n13 0.025
R1230 vss.n30 vss.n29 9.3
R1231 vss.n28 vss.n27 9.3
R1232 vss.n25 vss.n24 9.3
R1233 vss.n23 vss.n22 9.3
R1234 vss.n20 vss.n19 9.3
R1235 vss.n18 vss.n17 9.3
R1236 vss.n15 vss.n14 9.3
R1237 vss.n13 vss.n12 9.3
R1238 vss.n10 vss.n9 9.3
R1239 vss.n8 vss.n7 9.3
R1240 vss.n5 vss.n4 9.3
R1241 vss.n63 vss.n62 9.3
R1242 vss.n61 vss.n60 9.3
R1243 vss.n58 vss.n57 9.3
R1244 vss.n56 vss.n55 9.3
R1245 vss.n53 vss.n52 9.3
R1246 vss.n51 vss.n50 9.3
R1247 vss.n48 vss.n47 9.3
R1248 vss.n46 vss.n45 9.3
R1249 vss.n43 vss.n42 9.3
R1250 vss.n41 vss.n40 9.3
R1251 vss.n38 vss.n37 9.3
R1252 vss.n97 vss.n96 9.3
R1253 vss.n95 vss.n94 9.3
R1254 vss.n92 vss.n91 9.3
R1255 vss.n90 vss.n89 9.3
R1256 vss.n87 vss.n86 9.3
R1257 vss.n85 vss.n84 9.3
R1258 vss.n82 vss.n81 9.3
R1259 vss.n80 vss.n79 9.3
R1260 vss.n77 vss.n76 9.3
R1261 vss.n75 vss.n74 9.3
R1262 vss.n72 vss.n71 9.3
R1263 vss.n131 vss.n130 9.3
R1264 vss.n129 vss.n128 9.3
R1265 vss.n126 vss.n125 9.3
R1266 vss.n124 vss.n123 9.3
R1267 vss.n121 vss.n120 9.3
R1268 vss.n119 vss.n118 9.3
R1269 vss.n116 vss.n115 9.3
R1270 vss.n114 vss.n113 9.3
R1271 vss.n111 vss.n110 9.3
R1272 vss.n109 vss.n108 9.3
R1273 vss.n106 vss.n105 9.3
R1274 vss.n165 vss.n164 9.3
R1275 vss.n163 vss.n162 9.3
R1276 vss.n160 vss.n159 9.3
R1277 vss.n158 vss.n157 9.3
R1278 vss.n155 vss.n154 9.3
R1279 vss.n153 vss.n152 9.3
R1280 vss.n150 vss.n149 9.3
R1281 vss.n148 vss.n147 9.3
R1282 vss.n145 vss.n144 9.3
R1283 vss.n143 vss.n142 9.3
R1284 vss.n140 vss.n139 9.3
R1285 vss.n199 vss.n198 9.3
R1286 vss.n197 vss.n196 9.3
R1287 vss.n194 vss.n193 9.3
R1288 vss.n192 vss.n191 9.3
R1289 vss.n189 vss.n188 9.3
R1290 vss.n187 vss.n186 9.3
R1291 vss.n184 vss.n183 9.3
R1292 vss.n182 vss.n181 9.3
R1293 vss.n179 vss.n178 9.3
R1294 vss.n177 vss.n176 9.3
R1295 vss.n174 vss.n173 9.3
R1296 vss.n233 vss.n232 9.3
R1297 vss.n231 vss.n230 9.3
R1298 vss.n228 vss.n227 9.3
R1299 vss.n226 vss.n225 9.3
R1300 vss.n223 vss.n222 9.3
R1301 vss.n221 vss.n220 9.3
R1302 vss.n218 vss.n217 9.3
R1303 vss.n216 vss.n215 9.3
R1304 vss.n213 vss.n212 9.3
R1305 vss.n211 vss.n210 9.3
R1306 vss.n208 vss.n207 9.3
R1307 vss.n27 vss.n26 9.154
R1308 vss.n22 vss.n21 9.154
R1309 vss.n17 vss.n16 9.154
R1310 vss.n12 vss.n11 9.154
R1311 vss.n7 vss.n6 9.154
R1312 vss.n1 vss.n0 9.154
R1313 vss.n60 vss.n59 9.154
R1314 vss.n55 vss.n54 9.154
R1315 vss.n50 vss.n49 9.154
R1316 vss.n45 vss.n44 9.154
R1317 vss.n40 vss.n39 9.154
R1318 vss.n34 vss.n33 9.154
R1319 vss.n94 vss.n93 9.154
R1320 vss.n89 vss.n88 9.154
R1321 vss.n84 vss.n83 9.154
R1322 vss.n79 vss.n78 9.154
R1323 vss.n74 vss.n73 9.154
R1324 vss.n68 vss.n67 9.154
R1325 vss.n128 vss.n127 9.154
R1326 vss.n123 vss.n122 9.154
R1327 vss.n118 vss.n117 9.154
R1328 vss.n113 vss.n112 9.154
R1329 vss.n108 vss.n107 9.154
R1330 vss.n102 vss.n101 9.154
R1331 vss.n162 vss.n161 9.154
R1332 vss.n157 vss.n156 9.154
R1333 vss.n152 vss.n151 9.154
R1334 vss.n147 vss.n146 9.154
R1335 vss.n142 vss.n141 9.154
R1336 vss.n136 vss.n135 9.154
R1337 vss.n196 vss.n195 9.154
R1338 vss.n191 vss.n190 9.154
R1339 vss.n186 vss.n185 9.154
R1340 vss.n181 vss.n180 9.154
R1341 vss.n176 vss.n175 9.154
R1342 vss.n170 vss.n169 9.154
R1343 vss.n230 vss.n229 9.154
R1344 vss.n225 vss.n224 9.154
R1345 vss.n220 vss.n219 9.154
R1346 vss.n215 vss.n214 9.154
R1347 vss.n210 vss.n209 9.154
R1348 vss.n204 vss.n203 9.154
R1349 vss.n235 vss.n234 6.208
R1350 vss.n206 vss.n204 5.875
R1351 vss.n65 vss.n64 5.64
R1352 vss.n99 vss.n98 5.64
R1353 vss.n133 vss.n132 5.64
R1354 vss.n167 vss.n166 5.64
R1355 vss.n201 vss.n200 5.64
R1356 vss.n32 vss.n31 5.638
R1357 vss.n238 vss.n237 5.378
R1358 vss.n36 vss.n34 4.27
R1359 vss.n70 vss.n68 4.27
R1360 vss.n104 vss.n102 4.27
R1361 vss.n138 vss.n136 4.27
R1362 vss.n172 vss.n170 4.27
R1363 vss.n3 vss.n1 4.269
R1364 vss.n2 vss.t1 3.48
R1365 vss.n35 vss.t3 3.48
R1366 vss.n35 vss.t7 3.48
R1367 vss.n69 vss.t13 3.48
R1368 vss.n69 vss.t2 3.48
R1369 vss.n103 vss.t6 3.48
R1370 vss.n103 vss.t10 3.48
R1371 vss.n137 vss.t11 3.48
R1372 vss.n137 vss.t4 3.48
R1373 vss.n171 vss.t5 3.48
R1374 vss.n171 vss.t12 3.48
R1375 vss.n205 vss.t0 3.48
R1376 vss.n238 vss.n236 0.707
R1377 vss.n66 vss.n32 0.65
R1378 vss.n100 vss.n66 0.437
R1379 vss.n134 vss.n100 0.437
R1380 vss.n168 vss.n134 0.437
R1381 vss.n202 vss.n168 0.437
R1382 vss.n236 vss.n202 0.433
R1383 vss.n237 vss.t8 0.362
R1384 vss.n66 vss.n65 0.207
R1385 vss.n100 vss.n99 0.207
R1386 vss.n134 vss.n133 0.207
R1387 vss.n168 vss.n167 0.207
R1388 vss.n202 vss.n201 0.207
R1389 vss.n236 vss.n235 0.201
R1390 vss.n237 vss.t9 0.153
R1391 vss.n32 vss.n30 0.041
R1392 vss.n208 vss.n206 0.04
R1393 vss.n5 vss.n3 0.038
R1394 vss.n235 vss.n233 0.034
R1395 vss.n65 vss.n63 0.031
R1396 vss.n99 vss.n97 0.031
R1397 vss.n133 vss.n131 0.031
R1398 vss.n167 vss.n165 0.031
R1399 vss.n201 vss.n199 0.031
R1400 vss.n38 vss.n36 0.029
R1401 vss.n72 vss.n70 0.029
R1402 vss.n106 vss.n104 0.029
R1403 vss.n140 vss.n138 0.029
R1404 vss.n174 vss.n172 0.029
R1405 vss.n8 vss.n5 0.028
R1406 vss.n10 vss.n8 0.028
R1407 vss.n13 vss.n10 0.028
R1408 vss.n15 vss.n13 0.028
R1409 vss.n18 vss.n15 0.028
R1410 vss.n20 vss.n18 0.028
R1411 vss.n23 vss.n20 0.028
R1412 vss.n25 vss.n23 0.028
R1413 vss.n28 vss.n25 0.028
R1414 vss.n30 vss.n28 0.028
R1415 vss.n211 vss.n208 0.027
R1416 vss.n213 vss.n211 0.027
R1417 vss.n216 vss.n213 0.027
R1418 vss.n218 vss.n216 0.027
R1419 vss.n221 vss.n218 0.027
R1420 vss.n223 vss.n221 0.027
R1421 vss.n226 vss.n223 0.027
R1422 vss.n228 vss.n226 0.027
R1423 vss.n231 vss.n228 0.027
R1424 vss.n233 vss.n231 0.027
R1425 vss vss.n238 0.027
R1426 vss.n206 vss.n205 0.026
R1427 vss.n41 vss.n38 0.021
R1428 vss.n43 vss.n41 0.021
R1429 vss.n46 vss.n43 0.021
R1430 vss.n48 vss.n46 0.021
R1431 vss.n51 vss.n48 0.021
R1432 vss.n53 vss.n51 0.021
R1433 vss.n56 vss.n53 0.021
R1434 vss.n58 vss.n56 0.021
R1435 vss.n61 vss.n58 0.021
R1436 vss.n63 vss.n61 0.021
R1437 vss.n75 vss.n72 0.021
R1438 vss.n77 vss.n75 0.021
R1439 vss.n80 vss.n77 0.021
R1440 vss.n82 vss.n80 0.021
R1441 vss.n85 vss.n82 0.021
R1442 vss.n87 vss.n85 0.021
R1443 vss.n90 vss.n87 0.021
R1444 vss.n92 vss.n90 0.021
R1445 vss.n95 vss.n92 0.021
R1446 vss.n97 vss.n95 0.021
R1447 vss.n109 vss.n106 0.021
R1448 vss.n111 vss.n109 0.021
R1449 vss.n114 vss.n111 0.021
R1450 vss.n116 vss.n114 0.021
R1451 vss.n119 vss.n116 0.021
R1452 vss.n121 vss.n119 0.021
R1453 vss.n124 vss.n121 0.021
R1454 vss.n126 vss.n124 0.021
R1455 vss.n129 vss.n126 0.021
R1456 vss.n131 vss.n129 0.021
R1457 vss.n143 vss.n140 0.021
R1458 vss.n145 vss.n143 0.021
R1459 vss.n148 vss.n145 0.021
R1460 vss.n150 vss.n148 0.021
R1461 vss.n153 vss.n150 0.021
R1462 vss.n155 vss.n153 0.021
R1463 vss.n158 vss.n155 0.021
R1464 vss.n160 vss.n158 0.021
R1465 vss.n163 vss.n160 0.021
R1466 vss.n165 vss.n163 0.021
R1467 vss.n177 vss.n174 0.021
R1468 vss.n179 vss.n177 0.021
R1469 vss.n182 vss.n179 0.021
R1470 vss.n184 vss.n182 0.021
R1471 vss.n187 vss.n184 0.021
R1472 vss.n189 vss.n187 0.021
R1473 vss.n192 vss.n189 0.021
R1474 vss.n194 vss.n192 0.021
R1475 vss.n197 vss.n194 0.021
R1476 vss.n199 vss.n197 0.021
R1477 vss.n3 vss.n2 0.008
R1478 vss.n36 vss.n35 0.006
R1479 vss.n70 vss.n69 0.006
R1480 vss.n104 vss.n103 0.006
R1481 vss.n138 vss.n137 0.006
R1482 vss.n172 vss.n171 0.006
R1483 vinp.n14 vinp.t18 354.042
R1484 vinp.n16 vinp.t21 354.034
R1485 vinp.n20 vinp.t20 354.033
R1486 vinp.n20 vinp.t22 354.033
R1487 vinp.n16 vinp.t17 354.031
R1488 vinp.n14 vinp.t15 354.025
R1489 vinp.n13 vinp.t14 194.319
R1490 vinp.n21 vinp.t16 194.297
R1491 vinp.n21 vinp.t24 194.297
R1492 vinp.n17 vinp.t13 194.297
R1493 vinp.n17 vinp.t25 194.297
R1494 vinp.n13 vinp.t23 194.294
R1495 vinp.n22 vinp.n20 179.283
R1496 vinp.n15 vinp.n14 179.276
R1497 vinp.n18 vinp.n16 179.189
R1498 vinp.n15 vinp.n13 97.45
R1499 vinp.n22 vinp.n21 97.396
R1500 vinp.n18 vinp.n17 97.268
R1501 vinp.n28 vinp.t2 5.713
R1502 vinp.n28 vinp.t0 5.713
R1503 vinp.n26 vinp.t8 5.713
R1504 vinp.n26 vinp.t1 5.713
R1505 vinp.n32 vinp.t11 5.713
R1506 vinp.n32 vinp.t5 5.713
R1507 vinp.n27 vinp.t9 3.48
R1508 vinp.n27 vinp.t3 3.48
R1509 vinp.n25 vinp.t10 3.48
R1510 vinp.n25 vinp.t7 3.48
R1511 vinp.n31 vinp.t6 3.48
R1512 vinp.n31 vinp.t4 3.48
R1513 vinp.n24 vinp.n23 2.751
R1514 vinp.n1 vinp 1.25
R1515 vinp.n0 vinp 1.162
R1516 vinp.n4 vinp 0.973
R1517 vinp.n3 vinp 0.909
R1518 vinp.n23 vinp.n19 0.841
R1519 vinp.n19 vinp.n15 0.804
R1520 vinp.n7 vinp 0.696
R1521 vinp.n6 vinp 0.655
R1522 vinp.n10 vinp 0.418
R1523 vinp.n9 vinp 0.401
R1524 vinp.n26 vinp.n25 0.39
R1525 vinp.n32 vinp.n31 0.39
R1526 vinp.n28 vinp.n27 0.357
R1527 vinp.n33 vinp.n32 0.287
R1528 vinp.n29 vinp.n28 0.2
R1529 vinp.n30 vinp.n26 0.2
R1530 vinp.n30 vinp.n29 0.165
R1531 vinp.n12 vinp 0.147
R1532 vinp.n0 vinp.t19 0.14
R1533 vinp vinp.n34 0.139
R1534 vinp.n2 vinp.n1 0.117
R1535 vinp.n3 vinp.n2 0.117
R1536 vinp.n5 vinp.n4 0.117
R1537 vinp.n6 vinp.n5 0.117
R1538 vinp.n8 vinp.n7 0.117
R1539 vinp.n9 vinp.n8 0.117
R1540 vinp.n11 vinp.n10 0.117
R1541 vinp.n12 vinp.n11 0.117
R1542 vinp vinp.n33 0.096
R1543 vinp.n29 vinp.n24 0.076
R1544 vinp.n2 vinp.t12 0.023
R1545 vinp.n5 vinp.t27 0.023
R1546 vinp.n8 vinp.t28 0.023
R1547 vinp.n11 vinp.t26 0.023
R1548 vinp.n34 vinp.n12 0.021
R1549 vinp.n33 vinp.n30 0.02
R1550 vinp.n4 vinp.n3 0.019
R1551 vinp.n7 vinp.n6 0.019
R1552 vinp.n10 vinp.n9 0.019
R1553 vinp.n1 vinp.n0 0.018
R1554 vinp.n33 vinp.n24 0.011
R1555 vinp.n34 vinp 0.007
R1556 vinp.n19 vinp.n18 0.001
R1557 vinp.n23 vinp.n22 0.001
R1558 a_19910_7410.n7 a_19910_7410.t14 708.072
R1559 a_19910_7410.n9 a_19910_7410.t18 708.056
R1560 a_19910_7410.n11 a_19910_7410.t19 708.054
R1561 a_19910_7410.n11 a_19910_7410.t17 708.054
R1562 a_19910_7410.n9 a_19910_7410.t23 708.05
R1563 a_19910_7410.n7 a_19910_7410.t15 708.038
R1564 a_19910_7410.n6 a_19910_7410.t21 388.574
R1565 a_19910_7410.n6 a_19910_7410.t16 388.524
R1566 a_19910_7410.n12 a_19910_7410.t22 388.509
R1567 a_19910_7410.n12 a_19910_7410.t24 388.509
R1568 a_19910_7410.n10 a_19910_7410.t13 388.509
R1569 a_19910_7410.n10 a_19910_7410.t20 388.509
R1570 a_19910_7410.n13 a_19910_7410.t8 5.713
R1571 a_19910_7410.n13 a_19910_7410.t2 5.713
R1572 a_19910_7410.n5 a_19910_7410.t11 5.713
R1573 a_19910_7410.n5 a_19910_7410.t6 5.713
R1574 a_19910_7410.n3 a_19910_7410.t5 5.713
R1575 a_19910_7410.n3 a_19910_7410.t12 5.713
R1576 a_19910_7410.n4 a_19910_7410.t1 3.48
R1577 a_19910_7410.n4 a_19910_7410.t3 3.48
R1578 a_19910_7410.n2 a_19910_7410.t4 3.48
R1579 a_19910_7410.n2 a_19910_7410.t7 3.48
R1580 a_19910_7410.t0 a_19910_7410.n14 3.48
R1581 a_19910_7410.n14 a_19910_7410.t9 3.48
R1582 a_19910_7410.t10 a_19910_7410.n1 2.751
R1583 a_19910_7410.n1 a_19910_7410.n11 2.272
R1584 a_19910_7410.n8 a_19910_7410.n7 2.265
R1585 a_19910_7410.n0 a_19910_7410.n9 2.178
R1586 a_19910_7410.n14 a_19910_7410.n13 1.165
R1587 a_19910_7410.n5 a_19910_7410.n4 1.164
R1588 a_19910_7410.n3 a_19910_7410.n2 1.111
R1589 a_19910_7410.n1 a_19910_7410.n0 0.841
R1590 a_19910_7410.n0 a_19910_7410.n8 0.804
R1591 a_19910_7410.n8 a_19910_7410.n6 0.328
R1592 a_19910_7410.n1 a_19910_7410.n12 0.29
R1593 a_19910_7410.t10 a_19910_7410.n3 0.2
R1594 a_19910_7410.t10 a_19910_7410.n5 0.2
R1595 a_19910_7410.n13 a_19910_7410.t10 0.2
R1596 a_19910_7410.n0 a_19910_7410.n10 0.162
R1597 a_19840_7313.n7 a_19840_7313.t12 708.034
R1598 a_19840_7313.n6 a_19840_7313.t15 708.034
R1599 a_19840_7313.n9 a_19840_7313.t17 708.034
R1600 a_19840_7313.n7 a_19840_7313.t16 708.034
R1601 a_19840_7313.n6 a_19840_7313.t22 708.034
R1602 a_19840_7313.n9 a_19840_7313.t18 708.034
R1603 a_19840_7313.n10 a_19840_7313.t14 388.664
R1604 a_19840_7313.n8 a_19840_7313.t24 388.587
R1605 a_19840_7313.n8 a_19840_7313.t21 388.587
R1606 a_19840_7313.n5 a_19840_7313.t20 388.587
R1607 a_19840_7313.n5 a_19840_7313.t13 388.587
R1608 a_19840_7313.n10 a_19840_7313.t19 388.543
R1609 a_19840_7313.n18 a_19840_7313.t0 5.713
R1610 a_19840_7313.n18 a_19840_7313.t1 5.713
R1611 a_19840_7313.n14 a_19840_7313.t2 5.713
R1612 a_19840_7313.n14 a_19840_7313.t3 5.713
R1613 a_19840_7313.n3 a_19840_7313.t4 5.713
R1614 a_19840_7313.n3 a_19840_7313.t11 5.713
R1615 a_19840_7313.n13 a_19840_7313.t5 3.48
R1616 a_19840_7313.n13 a_19840_7313.t7 3.48
R1617 a_19840_7313.n2 a_19840_7313.t6 3.48
R1618 a_19840_7313.n2 a_19840_7313.t8 3.48
R1619 a_19840_7313.n20 a_19840_7313.t9 3.48
R1620 a_19840_7313.t10 a_19840_7313.n20 3.48
R1621 a_19840_7313.n12 a_19840_7313.n0 2.556
R1622 a_19840_7313.n0 a_19840_7313.n6 2.489
R1623 a_19840_7313.n11 a_19840_7313.n9 2.478
R1624 a_19840_7313.n1 a_19840_7313.n7 2.348
R1625 a_19840_7313.n0 a_19840_7313.n1 0.841
R1626 a_19840_7313.n1 a_19840_7313.n11 0.819
R1627 a_19840_7313.n15 a_19840_7313.n13 0.701
R1628 a_19840_7313.n4 a_19840_7313.n2 0.701
R1629 a_19840_7313.n20 a_19840_7313.n19 0.701
R1630 a_19840_7313.n15 a_19840_7313.n14 0.463
R1631 a_19840_7313.n4 a_19840_7313.n3 0.463
R1632 a_19840_7313.n19 a_19840_7313.n18 0.419
R1633 a_19840_7313.t23 a_19840_7313.n4 0.141
R1634 a_19840_7313.n17 a_19840_7313.n16 0.135
R1635 a_19840_7313.n16 a_19840_7313.n15 0.116
R1636 a_19840_7313.n19 a_19840_7313.n17 0.112
R1637 a_19840_7313.n11 a_19840_7313.n10 0.099
R1638 a_19840_7313.n0 a_19840_7313.n5 0.077
R1639 a_19840_7313.n17 a_19840_7313.n12 0.058
R1640 a_19840_7313.n1 a_19840_7313.n8 0.03
R1641 a_19840_7313.n12 a_19840_7313.t23 0.025
R1642 a_29168_7410.n4 a_29168_7410.t17 708.072
R1643 a_29168_7410.n6 a_29168_7410.t19 708.056
R1644 a_29168_7410.n8 a_29168_7410.t21 708.054
R1645 a_29168_7410.n8 a_29168_7410.t16 708.054
R1646 a_29168_7410.n6 a_29168_7410.t20 708.05
R1647 a_29168_7410.n4 a_29168_7410.t23 708.038
R1648 a_29168_7410.n3 a_29168_7410.t24 388.574
R1649 a_29168_7410.n3 a_29168_7410.t18 388.524
R1650 a_29168_7410.n9 a_29168_7410.t22 388.509
R1651 a_29168_7410.n9 a_29168_7410.t13 388.509
R1652 a_29168_7410.n7 a_29168_7410.t14 388.509
R1653 a_29168_7410.n7 a_29168_7410.t15 388.509
R1654 a_29168_7410.n14 a_29168_7410.t7 5.713
R1655 a_29168_7410.n14 a_29168_7410.t2 5.713
R1656 a_29168_7410.n11 a_29168_7410.t1 5.713
R1657 a_29168_7410.n11 a_29168_7410.t9 5.713
R1658 a_29168_7410.n13 a_29168_7410.t0 5.713
R1659 a_29168_7410.n13 a_29168_7410.t12 5.713
R1660 a_29168_7410.n10 a_29168_7410.t11 3.48
R1661 a_29168_7410.n10 a_29168_7410.t5 3.48
R1662 a_29168_7410.n12 a_29168_7410.t4 3.48
R1663 a_29168_7410.n12 a_29168_7410.t6 3.48
R1664 a_29168_7410.t3 a_29168_7410.n15 3.48
R1665 a_29168_7410.n15 a_29168_7410.t8 3.48
R1666 a_29168_7410.n0 a_29168_7410.n2 2.751
R1667 a_29168_7410.n2 a_29168_7410.n8 2.272
R1668 a_29168_7410.n5 a_29168_7410.n4 2.265
R1669 a_29168_7410.n1 a_29168_7410.n6 2.178
R1670 a_29168_7410.n11 a_29168_7410.n10 1.164
R1671 a_29168_7410.n13 a_29168_7410.n12 1.164
R1672 a_29168_7410.n15 a_29168_7410.n14 1.112
R1673 a_29168_7410.n2 a_29168_7410.n1 0.841
R1674 a_29168_7410.n1 a_29168_7410.n5 0.804
R1675 a_29168_7410.n0 a_29168_7410.n13 0.342
R1676 a_29168_7410.n5 a_29168_7410.n3 0.328
R1677 a_29168_7410.n2 a_29168_7410.n9 0.29
R1678 a_29168_7410.n0 a_29168_7410.n11 0.2
R1679 a_29168_7410.n14 a_29168_7410.n0 0.2
R1680 a_29168_7410.n1 a_29168_7410.n7 0.162
R1681 a_29168_7410.n0 a_29168_7410.t10 0.049
R1682 a_29098_7313.n7 a_29098_7313.t16 708.034
R1683 a_29098_7313.n6 a_29098_7313.t15 708.034
R1684 a_29098_7313.n8 a_29098_7313.t17 708.034
R1685 a_29098_7313.n7 a_29098_7313.t22 708.034
R1686 a_29098_7313.n6 a_29098_7313.t19 708.034
R1687 a_29098_7313.n8 a_29098_7313.t24 708.034
R1688 a_29098_7313.n9 a_29098_7313.t20 388.664
R1689 a_29098_7313.n0 a_29098_7313.t14 388.587
R1690 a_29098_7313.n0 a_29098_7313.t21 388.587
R1691 a_29098_7313.n5 a_29098_7313.t18 388.587
R1692 a_29098_7313.n5 a_29098_7313.t13 388.587
R1693 a_29098_7313.n9 a_29098_7313.t23 388.543
R1694 a_29098_7313.n18 a_29098_7313.t7 5.713
R1695 a_29098_7313.n18 a_29098_7313.t8 5.713
R1696 a_29098_7313.n3 a_29098_7313.t1 5.713
R1697 a_29098_7313.n3 a_29098_7313.t3 5.713
R1698 a_29098_7313.n14 a_29098_7313.t11 5.713
R1699 a_29098_7313.n14 a_29098_7313.t0 5.713
R1700 a_29098_7313.n2 a_29098_7313.t10 3.48
R1701 a_29098_7313.n2 a_29098_7313.t6 3.48
R1702 a_29098_7313.n13 a_29098_7313.t5 3.48
R1703 a_29098_7313.n13 a_29098_7313.t4 3.48
R1704 a_29098_7313.n20 a_29098_7313.t9 3.48
R1705 a_29098_7313.t2 a_29098_7313.n20 3.48
R1706 a_29098_7313.n11 a_29098_7313.n1 2.556
R1707 a_29098_7313.n1 a_29098_7313.n6 2.489
R1708 a_29098_7313.n10 a_29098_7313.n8 2.478
R1709 a_29098_7313.n0 a_29098_7313.n7 2.348
R1710 a_29098_7313.n0 a_29098_7313.n10 0.848
R1711 a_29098_7313.n1 a_29098_7313.n0 0.841
R1712 a_29098_7313.n4 a_29098_7313.n2 0.701
R1713 a_29098_7313.n15 a_29098_7313.n13 0.701
R1714 a_29098_7313.n20 a_29098_7313.n19 0.701
R1715 a_29098_7313.n15 a_29098_7313.n14 0.463
R1716 a_29098_7313.n19 a_29098_7313.n18 0.463
R1717 a_29098_7313.n4 a_29098_7313.n3 0.419
R1718 a_29098_7313.n16 a_29098_7313.t12 0.388
R1719 a_29098_7313.n17 a_29098_7313.n16 0.148
R1720 a_29098_7313.n17 a_29098_7313.n12 0.135
R1721 a_29098_7313.n16 a_29098_7313.n15 0.116
R1722 a_29098_7313.n19 a_29098_7313.n17 0.116
R1723 a_29098_7313.n12 a_29098_7313.n4 0.112
R1724 a_29098_7313.n10 a_29098_7313.n9 0.099
R1725 a_29098_7313.n1 a_29098_7313.n5 0.077
R1726 a_29098_7313.n12 a_29098_7313.n11 0.058
R1727 vrec.n329 vrec.t12 112.822
R1728 vrec.n373 vrec.t16 112.822
R1729 vrec.n373 vrec.t6 112.822
R1730 vrec.n480 vrec.t10 112.822
R1731 vrec.n480 vrec.t18 112.822
R1732 vrec.n6 vrec.t20 112.822
R1733 vrec.n6 vrec.t8 112.822
R1734 vrec.n71 vrec.t2 112.822
R1735 vrec.n71 vrec.t22 112.822
R1736 vrec.n252 vrec.t14 112.822
R1737 vrec.n252 vrec.t0 112.822
R1738 vrec.n147 vrec.t4 112.822
R1739 vrec.n13 vrec.n10 20.092
R1740 vrec.n297 vrec.n296 16.607
R1741 vrec.n220 vrec.n219 16.289
R1742 vrec.n70 vrec.n69 16.289
R1743 vrec.n448 vrec.n447 16.289
R1744 vrec.n372 vrec.n371 16.289
R1745 vrec.n155 vrec.n151 12.923
R1746 vrec.n302 vrec.n298 12.641
R1747 vrec.n381 vrec.n377 12.629
R1748 vrec.n453 vrec.n449 12.629
R1749 vrec.n79 vrec.n75 12.629
R1750 vrec.n225 vrec.n221 12.629
R1751 vrec.n145 vrec.n144 12.369
R1752 vrec.n304 vrec.n303 9.3
R1753 vrec.n310 vrec.n309 9.3
R1754 vrec.n316 vrec.n315 9.3
R1755 vrec.n322 vrec.n321 9.3
R1756 vrec.n328 vrec.n327 9.3
R1757 vrec.n340 vrec.n339 9.3
R1758 vrec.n346 vrec.n345 9.3
R1759 vrec.n352 vrec.n351 9.3
R1760 vrec.n358 vrec.n357 9.3
R1761 vrec.n364 vrec.n363 9.3
R1762 vrec.n369 vrec.n368 9.3
R1763 vrec.n383 vrec.n382 9.3
R1764 vrec.n389 vrec.n388 9.3
R1765 vrec.n395 vrec.n394 9.3
R1766 vrec.n401 vrec.n400 9.3
R1767 vrec.n407 vrec.n406 9.3
R1768 vrec.n415 vrec.n414 9.3
R1769 vrec.n421 vrec.n420 9.3
R1770 vrec.n427 vrec.n426 9.3
R1771 vrec.n433 vrec.n432 9.3
R1772 vrec.n439 vrec.n438 9.3
R1773 vrec.n444 vrec.n443 9.3
R1774 vrec.n455 vrec.n454 9.3
R1775 vrec.n461 vrec.n460 9.3
R1776 vrec.n467 vrec.n466 9.3
R1777 vrec.n473 vrec.n472 9.3
R1778 vrec.n479 vrec.n478 9.3
R1779 vrec.n491 vrec.n490 9.3
R1780 vrec.n497 vrec.n496 9.3
R1781 vrec.n503 vrec.n502 9.3
R1782 vrec.n509 vrec.n508 9.3
R1783 vrec.n515 vrec.n514 9.3
R1784 vrec.n520 vrec.n519 9.3
R1785 vrec.n81 vrec.n80 9.3
R1786 vrec.n87 vrec.n86 9.3
R1787 vrec.n93 vrec.n92 9.3
R1788 vrec.n99 vrec.n98 9.3
R1789 vrec.n105 vrec.n104 9.3
R1790 vrec.n113 vrec.n112 9.3
R1791 vrec.n119 vrec.n118 9.3
R1792 vrec.n125 vrec.n124 9.3
R1793 vrec.n131 vrec.n130 9.3
R1794 vrec.n137 vrec.n136 9.3
R1795 vrec.n142 vrec.n141 9.3
R1796 vrec.n217 vrec.n216 9.3
R1797 vrec.n157 vrec.n156 9.3
R1798 vrec.n163 vrec.n162 9.3
R1799 vrec.n169 vrec.n168 9.3
R1800 vrec.n175 vrec.n174 9.3
R1801 vrec.n181 vrec.n180 9.3
R1802 vrec.n189 vrec.n188 9.3
R1803 vrec.n195 vrec.n194 9.3
R1804 vrec.n201 vrec.n200 9.3
R1805 vrec.n207 vrec.n206 9.3
R1806 vrec.n212 vrec.n211 9.3
R1807 vrec.n227 vrec.n226 9.3
R1808 vrec.n233 vrec.n232 9.3
R1809 vrec.n239 vrec.n238 9.3
R1810 vrec.n245 vrec.n244 9.3
R1811 vrec.n251 vrec.n250 9.3
R1812 vrec.n263 vrec.n262 9.3
R1813 vrec.n269 vrec.n268 9.3
R1814 vrec.n275 vrec.n274 9.3
R1815 vrec.n281 vrec.n280 9.3
R1816 vrec.n287 vrec.n286 9.3
R1817 vrec.n292 vrec.n291 9.3
R1818 vrec.n231 vrec.n230 9.3
R1819 vrec.n237 vrec.n236 9.3
R1820 vrec.n243 vrec.n242 9.3
R1821 vrec.n249 vrec.n248 9.3
R1822 vrec.n267 vrec.n266 9.3
R1823 vrec.n273 vrec.n272 9.3
R1824 vrec.n279 vrec.n278 9.3
R1825 vrec.n285 vrec.n284 9.3
R1826 vrec.n290 vrec.n289 9.3
R1827 vrec.n85 vrec.n84 9.3
R1828 vrec.n91 vrec.n90 9.3
R1829 vrec.n97 vrec.n96 9.3
R1830 vrec.n103 vrec.n102 9.3
R1831 vrec.n117 vrec.n116 9.3
R1832 vrec.n123 vrec.n122 9.3
R1833 vrec.n129 vrec.n128 9.3
R1834 vrec.n135 vrec.n134 9.3
R1835 vrec.n140 vrec.n139 9.3
R1836 vrec.n459 vrec.n458 9.3
R1837 vrec.n465 vrec.n464 9.3
R1838 vrec.n471 vrec.n470 9.3
R1839 vrec.n477 vrec.n476 9.3
R1840 vrec.n495 vrec.n494 9.3
R1841 vrec.n501 vrec.n500 9.3
R1842 vrec.n507 vrec.n506 9.3
R1843 vrec.n513 vrec.n512 9.3
R1844 vrec.n518 vrec.n517 9.3
R1845 vrec.n387 vrec.n386 9.3
R1846 vrec.n393 vrec.n392 9.3
R1847 vrec.n399 vrec.n398 9.3
R1848 vrec.n405 vrec.n404 9.3
R1849 vrec.n419 vrec.n418 9.3
R1850 vrec.n425 vrec.n424 9.3
R1851 vrec.n431 vrec.n430 9.3
R1852 vrec.n437 vrec.n436 9.3
R1853 vrec.n442 vrec.n441 9.3
R1854 vrec.n308 vrec.n307 9.3
R1855 vrec.n314 vrec.n313 9.3
R1856 vrec.n320 vrec.n319 9.3
R1857 vrec.n326 vrec.n325 9.3
R1858 vrec.n344 vrec.n343 9.3
R1859 vrec.n350 vrec.n349 9.3
R1860 vrec.n356 vrec.n355 9.3
R1861 vrec.n362 vrec.n361 9.3
R1862 vrec.n367 vrec.n366 9.3
R1863 vrec.n161 vrec.n160 9.3
R1864 vrec.n167 vrec.n166 9.3
R1865 vrec.n173 vrec.n172 9.3
R1866 vrec.n179 vrec.n178 9.3
R1867 vrec.n193 vrec.n192 9.3
R1868 vrec.n199 vrec.n198 9.3
R1869 vrec.n205 vrec.n204 9.3
R1870 vrec.n210 vrec.n209 9.3
R1871 vrec.n215 vrec.n214 9.3
R1872 vrec.n15 vrec.n14 9.3
R1873 vrec.n18 vrec.n17 9.3
R1874 vrec.n20 vrec.n19 9.3
R1875 vrec.n23 vrec.n22 9.3
R1876 vrec.n25 vrec.n24 9.3
R1877 vrec.n28 vrec.n27 9.3
R1878 vrec.n30 vrec.n29 9.3
R1879 vrec.n33 vrec.n32 9.3
R1880 vrec.n35 vrec.n34 9.3
R1881 vrec.n42 vrec.n41 9.3
R1882 vrec.n45 vrec.n44 9.3
R1883 vrec.n47 vrec.n46 9.3
R1884 vrec.n50 vrec.n49 9.3
R1885 vrec.n52 vrec.n51 9.3
R1886 vrec.n55 vrec.n54 9.3
R1887 vrec.n57 vrec.n56 9.3
R1888 vrec.n60 vrec.n59 9.3
R1889 vrec.n62 vrec.n61 9.3
R1890 vrec.n65 vrec.n64 9.3
R1891 vrec.n67 vrec.n66 9.3
R1892 vrec.n224 vrec.n223 8.855
R1893 vrec.n230 vrec.n229 8.855
R1894 vrec.n236 vrec.n235 8.855
R1895 vrec.n242 vrec.n241 8.855
R1896 vrec.n248 vrec.n247 8.855
R1897 vrec.n255 vrec.n254 8.855
R1898 vrec.n260 vrec.n259 8.855
R1899 vrec.n266 vrec.n265 8.855
R1900 vrec.n272 vrec.n271 8.855
R1901 vrec.n278 vrec.n277 8.855
R1902 vrec.n284 vrec.n283 8.855
R1903 vrec.n289 vrec.n288 8.855
R1904 vrec.n78 vrec.n77 8.855
R1905 vrec.n84 vrec.n83 8.855
R1906 vrec.n90 vrec.n89 8.855
R1907 vrec.n96 vrec.n95 8.855
R1908 vrec.n102 vrec.n101 8.855
R1909 vrec.n74 vrec.n73 8.855
R1910 vrec.n110 vrec.n109 8.855
R1911 vrec.n116 vrec.n115 8.855
R1912 vrec.n122 vrec.n121 8.855
R1913 vrec.n128 vrec.n127 8.855
R1914 vrec.n134 vrec.n133 8.855
R1915 vrec.n139 vrec.n138 8.855
R1916 vrec.n452 vrec.n451 8.855
R1917 vrec.n458 vrec.n457 8.855
R1918 vrec.n464 vrec.n463 8.855
R1919 vrec.n470 vrec.n469 8.855
R1920 vrec.n476 vrec.n475 8.855
R1921 vrec.n483 vrec.n482 8.855
R1922 vrec.n488 vrec.n487 8.855
R1923 vrec.n494 vrec.n493 8.855
R1924 vrec.n500 vrec.n499 8.855
R1925 vrec.n506 vrec.n505 8.855
R1926 vrec.n512 vrec.n511 8.855
R1927 vrec.n517 vrec.n516 8.855
R1928 vrec.n380 vrec.n379 8.855
R1929 vrec.n386 vrec.n385 8.855
R1930 vrec.n392 vrec.n391 8.855
R1931 vrec.n398 vrec.n397 8.855
R1932 vrec.n404 vrec.n403 8.855
R1933 vrec.n376 vrec.n375 8.855
R1934 vrec.n412 vrec.n411 8.855
R1935 vrec.n418 vrec.n417 8.855
R1936 vrec.n424 vrec.n423 8.855
R1937 vrec.n430 vrec.n429 8.855
R1938 vrec.n436 vrec.n435 8.855
R1939 vrec.n441 vrec.n440 8.855
R1940 vrec.n301 vrec.n300 8.855
R1941 vrec.n307 vrec.n306 8.855
R1942 vrec.n313 vrec.n312 8.855
R1943 vrec.n319 vrec.n318 8.855
R1944 vrec.n325 vrec.n324 8.855
R1945 vrec.n332 vrec.n331 8.855
R1946 vrec.n337 vrec.n336 8.855
R1947 vrec.n343 vrec.n342 8.855
R1948 vrec.n349 vrec.n348 8.855
R1949 vrec.n355 vrec.n354 8.855
R1950 vrec.n361 vrec.n360 8.855
R1951 vrec.n366 vrec.n365 8.855
R1952 vrec.n154 vrec.n153 8.855
R1953 vrec.n160 vrec.n159 8.855
R1954 vrec.n166 vrec.n165 8.855
R1955 vrec.n172 vrec.n171 8.855
R1956 vrec.n178 vrec.n177 8.855
R1957 vrec.n184 vrec.n183 8.855
R1958 vrec.n150 vrec.n149 8.855
R1959 vrec.n192 vrec.n191 8.855
R1960 vrec.n198 vrec.n197 8.855
R1961 vrec.n204 vrec.n203 8.855
R1962 vrec.n209 vrec.n208 8.855
R1963 vrec.n214 vrec.n213 8.855
R1964 vrec.n12 vrec.n11 8.855
R1965 vrec.n17 vrec.n16 8.855
R1966 vrec.n22 vrec.n21 8.855
R1967 vrec.n27 vrec.n26 8.855
R1968 vrec.n32 vrec.n31 8.855
R1969 vrec.n9 vrec.n8 8.855
R1970 vrec.n39 vrec.n38 8.855
R1971 vrec.n44 vrec.n43 8.855
R1972 vrec.n49 vrec.n48 8.855
R1973 vrec.n54 vrec.n53 8.855
R1974 vrec.n59 vrec.n58 8.855
R1975 vrec.n64 vrec.n63 8.855
R1976 vrec.n8 vrec.n7 7.463
R1977 vrec.n293 vrec.n220 6.209
R1978 vrec.n143 vrec.n70 6.209
R1979 vrec.n521 vrec.n448 6.209
R1980 vrec.n445 vrec.n372 6.209
R1981 vrec.n68 vrec.n0 6.209
R1982 vrec.n370 vrec.n297 6.208
R1983 vrec.n253 vrec.n252 5.95
R1984 vrec.n72 vrec.n71 5.95
R1985 vrec.n481 vrec.n480 5.95
R1986 vrec.n374 vrec.n373 5.95
R1987 vrec.n261 vrec.n260 5.876
R1988 vrec.n111 vrec.n110 5.876
R1989 vrec.n489 vrec.n488 5.876
R1990 vrec.n413 vrec.n412 5.876
R1991 vrec.n40 vrec.n39 5.876
R1992 vrec.n185 vrec.n184 5.873
R1993 vrec.n338 vrec.n337 5.873
R1994 vrec.n37 vrec.t21 5.713
R1995 vrec.n485 vrec.t11 5.713
R1996 vrec.n485 vrec.t19 5.713
R1997 vrec.n334 vrec.t13 5.713
R1998 vrec.n409 vrec.t17 5.713
R1999 vrec.n409 vrec.t7 5.713
R2000 vrec.n257 vrec.t15 5.713
R2001 vrec.n257 vrec.t1 5.713
R2002 vrec.n107 vrec.t3 5.713
R2003 vrec.n107 vrec.t23 5.713
R2004 vrec.n186 vrec.t5 5.713
R2005 vrec.n37 vrec.t9 5.713
R2006 vrec.n218 vrec.n145 5.637
R2007 vrec.n381 vrec.n380 5.614
R2008 vrec.n79 vrec.n78 5.614
R2009 vrec.n225 vrec.n224 5.614
R2010 vrec.n453 vrec.n452 5.614
R2011 vrec.n13 vrec.n12 5.614
R2012 vrec.n302 vrec.n301 5.611
R2013 vrec.n155 vrec.n154 5.571
R2014 vrec.n330 vrec.n329 5.347
R2015 vrec.n148 vrec.n147 5.347
R2016 vrec.n484 vrec.n483 4.27
R2017 vrec.n256 vrec.n255 4.27
R2018 vrec.n106 vrec.n74 4.27
R2019 vrec.n408 vrec.n376 4.27
R2020 vrec.n36 vrec.n9 4.27
R2021 vrec.n333 vrec.n332 4.269
R2022 vrec.n187 vrec.n150 4.269
R2023 vrec.n203 vrec.n202 3.685
R2024 vrec.n197 vrec.n196 3.685
R2025 vrec.n191 vrec.n190 3.685
R2026 vrec.n149 vrec.n148 3.685
R2027 vrec.n183 vrec.n182 3.685
R2028 vrec.n177 vrec.n176 3.685
R2029 vrec.n171 vrec.n170 3.685
R2030 vrec.n165 vrec.n164 3.685
R2031 vrec.n159 vrec.n158 3.685
R2032 vrec.n360 vrec.n359 3.685
R2033 vrec.n354 vrec.n353 3.685
R2034 vrec.n348 vrec.n347 3.685
R2035 vrec.n342 vrec.n341 3.685
R2036 vrec.n336 vrec.n335 3.685
R2037 vrec.n331 vrec.n330 3.685
R2038 vrec.n324 vrec.n323 3.685
R2039 vrec.n318 vrec.n317 3.685
R2040 vrec.n312 vrec.n311 3.685
R2041 vrec.n306 vrec.n305 3.685
R2042 vrec.n153 vrec.n152 3.514
R2043 vrec.n300 vrec.n299 3.514
R2044 vrec.n435 vrec.n434 3.052
R2045 vrec.n429 vrec.n428 3.052
R2046 vrec.n423 vrec.n422 3.052
R2047 vrec.n417 vrec.n416 3.052
R2048 vrec.n411 vrec.n410 3.052
R2049 vrec.n375 vrec.n374 3.052
R2050 vrec.n403 vrec.n402 3.052
R2051 vrec.n397 vrec.n396 3.052
R2052 vrec.n391 vrec.n390 3.052
R2053 vrec.n385 vrec.n384 3.052
R2054 vrec.n511 vrec.n510 3.052
R2055 vrec.n505 vrec.n504 3.052
R2056 vrec.n499 vrec.n498 3.052
R2057 vrec.n493 vrec.n492 3.052
R2058 vrec.n487 vrec.n486 3.052
R2059 vrec.n482 vrec.n481 3.052
R2060 vrec.n475 vrec.n474 3.052
R2061 vrec.n469 vrec.n468 3.052
R2062 vrec.n463 vrec.n462 3.052
R2063 vrec.n457 vrec.n456 3.052
R2064 vrec.n133 vrec.n132 3.052
R2065 vrec.n127 vrec.n126 3.052
R2066 vrec.n121 vrec.n120 3.052
R2067 vrec.n115 vrec.n114 3.052
R2068 vrec.n109 vrec.n108 3.052
R2069 vrec.n73 vrec.n72 3.052
R2070 vrec.n101 vrec.n100 3.052
R2071 vrec.n95 vrec.n94 3.052
R2072 vrec.n89 vrec.n88 3.052
R2073 vrec.n83 vrec.n82 3.052
R2074 vrec.n283 vrec.n282 3.052
R2075 vrec.n277 vrec.n276 3.052
R2076 vrec.n271 vrec.n270 3.052
R2077 vrec.n265 vrec.n264 3.052
R2078 vrec.n259 vrec.n258 3.052
R2079 vrec.n254 vrec.n253 3.052
R2080 vrec.n247 vrec.n246 3.052
R2081 vrec.n241 vrec.n240 3.052
R2082 vrec.n235 vrec.n234 3.052
R2083 vrec.n229 vrec.n228 3.052
R2084 vrec.n379 vrec.n378 2.91
R2085 vrec.n451 vrec.n450 2.91
R2086 vrec.n77 vrec.n76 2.91
R2087 vrec.n223 vrec.n222 2.91
R2088 vrec.n524 vrec.n523 2.18
R2089 vrec.n524 vrec.t25 0.868
R2090 vrec.n294 vrec.n218 0.768
R2091 vrec.n446 vrec.n370 0.75
R2092 vrec vrec.t24 0.749
R2093 vrec.n157 vrec.n155 0.713
R2094 vrec.n6 vrec.n5 0.697
R2095 vrec.n6 vrec.n4 0.697
R2096 vrec.n7 vrec.n6 0.697
R2097 vrec.n6 vrec.n3 0.697
R2098 vrec.n6 vrec.n2 0.697
R2099 vrec.n6 vrec.n1 0.697
R2100 vrec.n304 vrec.n302 0.668
R2101 vrec.n15 vrec.n13 0.652
R2102 vrec.n383 vrec.n381 0.652
R2103 vrec.n455 vrec.n453 0.652
R2104 vrec.n81 vrec.n79 0.652
R2105 vrec.n227 vrec.n225 0.652
R2106 vrec.n147 vrec.n146 0.592
R2107 vrec.n523 vrec.n522 0.57
R2108 vrec.n522 vrec.n446 0.57
R2109 vrec.n523 vrec.n295 0.57
R2110 vrec.n295 vrec.n294 0.57
R2111 vrec.n446 vrec.n445 0.208
R2112 vrec.n522 vrec.n521 0.208
R2113 vrec.n295 vrec.n143 0.208
R2114 vrec.n294 vrec.n293 0.208
R2115 vrec.n523 vrec.n68 0.208
R2116 vrec vrec.n524 0.06
R2117 vrec.n340 vrec.n338 0.047
R2118 vrec.n185 vrec.n181 0.046
R2119 vrec.n218 vrec.n217 0.045
R2120 vrec.n333 vrec.n328 0.043
R2121 vrec.n189 vrec.n187 0.042
R2122 vrec.n370 vrec.n369 0.04
R2123 vrec.n369 vrec.n367 0.032
R2124 vrec.n367 vrec.n364 0.032
R2125 vrec.n364 vrec.n362 0.032
R2126 vrec.n362 vrec.n358 0.032
R2127 vrec.n358 vrec.n356 0.032
R2128 vrec.n356 vrec.n352 0.032
R2129 vrec.n352 vrec.n350 0.032
R2130 vrec.n350 vrec.n346 0.032
R2131 vrec.n346 vrec.n344 0.032
R2132 vrec.n344 vrec.n340 0.032
R2133 vrec.n328 vrec.n326 0.032
R2134 vrec.n326 vrec.n322 0.032
R2135 vrec.n322 vrec.n320 0.032
R2136 vrec.n320 vrec.n316 0.032
R2137 vrec.n316 vrec.n314 0.032
R2138 vrec.n314 vrec.n310 0.032
R2139 vrec.n310 vrec.n308 0.032
R2140 vrec.n308 vrec.n304 0.032
R2141 vrec.n415 vrec.n413 0.031
R2142 vrec.n491 vrec.n489 0.031
R2143 vrec.n113 vrec.n111 0.031
R2144 vrec.n263 vrec.n261 0.031
R2145 vrec.n42 vrec.n40 0.031
R2146 vrec.n217 vrec.n215 0.031
R2147 vrec.n215 vrec.n212 0.031
R2148 vrec.n212 vrec.n210 0.031
R2149 vrec.n210 vrec.n207 0.031
R2150 vrec.n207 vrec.n205 0.031
R2151 vrec.n205 vrec.n201 0.031
R2152 vrec.n201 vrec.n199 0.031
R2153 vrec.n199 vrec.n195 0.031
R2154 vrec.n195 vrec.n193 0.031
R2155 vrec.n193 vrec.n189 0.031
R2156 vrec.n181 vrec.n179 0.031
R2157 vrec.n179 vrec.n175 0.031
R2158 vrec.n175 vrec.n173 0.031
R2159 vrec.n173 vrec.n169 0.031
R2160 vrec.n169 vrec.n167 0.031
R2161 vrec.n167 vrec.n163 0.031
R2162 vrec.n163 vrec.n161 0.031
R2163 vrec.n161 vrec.n157 0.031
R2164 vrec.n338 vrec.n334 0.031
R2165 vrec.n186 vrec.n185 0.03
R2166 vrec.n408 vrec.n407 0.029
R2167 vrec.n484 vrec.n479 0.029
R2168 vrec.n106 vrec.n105 0.029
R2169 vrec.n256 vrec.n251 0.029
R2170 vrec.n36 vrec.n35 0.029
R2171 vrec.n445 vrec.n444 0.027
R2172 vrec.n521 vrec.n520 0.027
R2173 vrec.n143 vrec.n142 0.027
R2174 vrec.n293 vrec.n292 0.027
R2175 vrec.n68 vrec.n67 0.027
R2176 vrec.n444 vrec.n442 0.021
R2177 vrec.n442 vrec.n439 0.021
R2178 vrec.n439 vrec.n437 0.021
R2179 vrec.n437 vrec.n433 0.021
R2180 vrec.n433 vrec.n431 0.021
R2181 vrec.n431 vrec.n427 0.021
R2182 vrec.n427 vrec.n425 0.021
R2183 vrec.n425 vrec.n421 0.021
R2184 vrec.n421 vrec.n419 0.021
R2185 vrec.n419 vrec.n415 0.021
R2186 vrec.n407 vrec.n405 0.021
R2187 vrec.n405 vrec.n401 0.021
R2188 vrec.n401 vrec.n399 0.021
R2189 vrec.n399 vrec.n395 0.021
R2190 vrec.n395 vrec.n393 0.021
R2191 vrec.n393 vrec.n389 0.021
R2192 vrec.n389 vrec.n387 0.021
R2193 vrec.n387 vrec.n383 0.021
R2194 vrec.n520 vrec.n518 0.021
R2195 vrec.n518 vrec.n515 0.021
R2196 vrec.n515 vrec.n513 0.021
R2197 vrec.n513 vrec.n509 0.021
R2198 vrec.n509 vrec.n507 0.021
R2199 vrec.n507 vrec.n503 0.021
R2200 vrec.n503 vrec.n501 0.021
R2201 vrec.n501 vrec.n497 0.021
R2202 vrec.n497 vrec.n495 0.021
R2203 vrec.n495 vrec.n491 0.021
R2204 vrec.n479 vrec.n477 0.021
R2205 vrec.n477 vrec.n473 0.021
R2206 vrec.n473 vrec.n471 0.021
R2207 vrec.n471 vrec.n467 0.021
R2208 vrec.n467 vrec.n465 0.021
R2209 vrec.n465 vrec.n461 0.021
R2210 vrec.n461 vrec.n459 0.021
R2211 vrec.n459 vrec.n455 0.021
R2212 vrec.n142 vrec.n140 0.021
R2213 vrec.n140 vrec.n137 0.021
R2214 vrec.n137 vrec.n135 0.021
R2215 vrec.n135 vrec.n131 0.021
R2216 vrec.n131 vrec.n129 0.021
R2217 vrec.n129 vrec.n125 0.021
R2218 vrec.n125 vrec.n123 0.021
R2219 vrec.n123 vrec.n119 0.021
R2220 vrec.n119 vrec.n117 0.021
R2221 vrec.n117 vrec.n113 0.021
R2222 vrec.n105 vrec.n103 0.021
R2223 vrec.n103 vrec.n99 0.021
R2224 vrec.n99 vrec.n97 0.021
R2225 vrec.n97 vrec.n93 0.021
R2226 vrec.n93 vrec.n91 0.021
R2227 vrec.n91 vrec.n87 0.021
R2228 vrec.n87 vrec.n85 0.021
R2229 vrec.n85 vrec.n81 0.021
R2230 vrec.n292 vrec.n290 0.021
R2231 vrec.n290 vrec.n287 0.021
R2232 vrec.n287 vrec.n285 0.021
R2233 vrec.n285 vrec.n281 0.021
R2234 vrec.n281 vrec.n279 0.021
R2235 vrec.n279 vrec.n275 0.021
R2236 vrec.n275 vrec.n273 0.021
R2237 vrec.n273 vrec.n269 0.021
R2238 vrec.n269 vrec.n267 0.021
R2239 vrec.n267 vrec.n263 0.021
R2240 vrec.n251 vrec.n249 0.021
R2241 vrec.n249 vrec.n245 0.021
R2242 vrec.n245 vrec.n243 0.021
R2243 vrec.n243 vrec.n239 0.021
R2244 vrec.n239 vrec.n237 0.021
R2245 vrec.n237 vrec.n233 0.021
R2246 vrec.n233 vrec.n231 0.021
R2247 vrec.n231 vrec.n227 0.021
R2248 vrec.n67 vrec.n65 0.021
R2249 vrec.n65 vrec.n62 0.021
R2250 vrec.n62 vrec.n60 0.021
R2251 vrec.n60 vrec.n57 0.021
R2252 vrec.n57 vrec.n55 0.021
R2253 vrec.n55 vrec.n52 0.021
R2254 vrec.n52 vrec.n50 0.021
R2255 vrec.n50 vrec.n47 0.021
R2256 vrec.n47 vrec.n45 0.021
R2257 vrec.n45 vrec.n42 0.021
R2258 vrec.n35 vrec.n33 0.021
R2259 vrec.n33 vrec.n30 0.021
R2260 vrec.n30 vrec.n28 0.021
R2261 vrec.n28 vrec.n25 0.021
R2262 vrec.n25 vrec.n23 0.021
R2263 vrec.n23 vrec.n20 0.021
R2264 vrec.n20 vrec.n18 0.021
R2265 vrec.n18 vrec.n15 0.021
R2266 vrec.n413 vrec.n409 0.021
R2267 vrec.n489 vrec.n485 0.021
R2268 vrec.n111 vrec.n107 0.021
R2269 vrec.n261 vrec.n257 0.021
R2270 vrec.n40 vrec.n37 0.021
R2271 vrec.n334 vrec.n333 0.009
R2272 vrec.n187 vrec.n186 0.009
R2273 vrec.n409 vrec.n408 0.006
R2274 vrec.n485 vrec.n484 0.006
R2275 vrec.n107 vrec.n106 0.006
R2276 vrec.n257 vrec.n256 0.006
R2277 vrec.n37 vrec.n36 0.006
R2278 vinn.n31 vinn.t25 354.028
R2279 vinn.n29 vinn.t23 354.028
R2280 vinn.n34 vinn.t26 354.028
R2281 vinn.n31 vinn.t19 354.028
R2282 vinn.n29 vinn.t21 354.028
R2283 vinn.n34 vinn.t20 354.028
R2284 vinn.n35 vinn.t27 194.35
R2285 vinn.n32 vinn.t28 194.316
R2286 vinn.n32 vinn.t18 194.316
R2287 vinn.n28 vinn.t24 194.316
R2288 vinn.n28 vinn.t17 194.316
R2289 vinn.n35 vinn.t22 194.29
R2290 vinn.n30 vinn.n29 179.493
R2291 vinn.n36 vinn.n34 179.482
R2292 vinn.n33 vinn.n31 179.352
R2293 vinn.n36 vinn.n35 97.241
R2294 vinn.n30 vinn.n28 97.212
R2295 vinn.n33 vinn.n32 97.165
R2296 vinn.n40 vinn.t9 5.713
R2297 vinn.n40 vinn.t7 5.713
R2298 vinn.n22 vinn.t5 5.713
R2299 vinn.n22 vinn.t10 5.713
R2300 vinn.n26 vinn.t8 5.713
R2301 vinn.n26 vinn.t6 5.713
R2302 vinn.n39 vinn.t16 3.48
R2303 vinn.n39 vinn.t14 3.48
R2304 vinn.n21 vinn.t15 3.48
R2305 vinn.n21 vinn.t12 3.48
R2306 vinn.n25 vinn.t13 3.48
R2307 vinn.n25 vinn.t11 3.48
R2308 vinn.n43 vinn.n38 2.555
R2309 vinn.n1 vinn 1.231
R2310 vinn.n0 vinn 1.139
R2311 vinn.n2 vinn 1.133
R2312 vinn.n6 vinn 0.981
R2313 vinn.n4 vinn 0.89
R2314 vinn.n5 vinn 0.89
R2315 vinn.n7 vinn 0.883
R2316 vinn.n38 vinn.n37 0.841
R2317 vinn.n37 vinn.n36 0.819
R2318 vinn.n11 vinn 0.703
R2319 vinn.n9 vinn 0.641
R2320 vinn.n10 vinn 0.64
R2321 vinn.n12 vinn 0.632
R2322 vinn.n16 vinn 0.426
R2323 vinn.n14 vinn 0.391
R2324 vinn.n15 vinn 0.389
R2325 vinn.n23 vinn.n22 0.384
R2326 vinn.n27 vinn.n26 0.384
R2327 vinn.n17 vinn 0.381
R2328 vinn.n41 vinn.n40 0.343
R2329 vinn.n44 vinn.n27 0.266
R2330 vinn.n24 vinn.n23 0.195
R2331 vinn.n42 vinn.n41 0.189
R2332 vinn.n0 vinn.t0 0.143
R2333 vinn.n19 vinn 0.142
R2334 vinn vinn.n45 0.139
R2335 vinn.n20 vinn 0.138
R2336 vinn.n3 vinn.n2 0.118
R2337 vinn.n4 vinn.n3 0.118
R2338 vinn.n8 vinn.n7 0.118
R2339 vinn.n9 vinn.n8 0.118
R2340 vinn.n13 vinn.n12 0.118
R2341 vinn.n14 vinn.n13 0.118
R2342 vinn.n18 vinn.n17 0.118
R2343 vinn.n19 vinn.n18 0.118
R2344 vinn.n45 vinn.n44 0.103
R2345 vinn.n43 vinn.n42 0.068
R2346 vinn.n44 vinn.n24 0.057
R2347 vinn.n18 vinn.t2 0.025
R2348 vinn.n13 vinn.t3 0.025
R2349 vinn.n8 vinn.t1 0.025
R2350 vinn.n3 vinn.t4 0.025
R2351 vinn.n45 vinn.n20 0.013
R2352 vinn.n44 vinn.n43 0.012
R2353 vinn.n1 vinn.n0 0.007
R2354 vinn.n45 vinn 0.007
R2355 vinn.n41 vinn.n39 0.006
R2356 vinn.n23 vinn.n21 0.006
R2357 vinn.n27 vinn.n25 0.006
R2358 vinn.n2 vinn.n1 0.004
R2359 vinn.n5 vinn.n4 0.004
R2360 vinn.n7 vinn.n6 0.004
R2361 vinn.n10 vinn.n9 0.004
R2362 vinn.n12 vinn.n11 0.004
R2363 vinn.n15 vinn.n14 0.004
R2364 vinn.n17 vinn.n16 0.004
R2365 vinn.n20 vinn.n19 0.004
R2366 vinn.n6 vinn.n5 0.003
R2367 vinn.n11 vinn.n10 0.003
R2368 vinn.n16 vinn.n15 0.003
R2369 vinn.n38 vinn.n30 0.001
R2370 vinn.n37 vinn.n33 0.001
R2371 w_570_7310.n456 w_570_7310.t31 112.822
R2372 w_570_7310.n0 w_570_7310.t23 112.822
R2373 w_570_7310.n0 w_570_7310.t16 112.822
R2374 w_570_7310.n359 w_570_7310.t6 112.822
R2375 w_570_7310.n359 w_570_7310.t33 112.822
R2376 w_570_7310.n52 w_570_7310.t27 112.822
R2377 w_570_7310.n52 w_570_7310.t8 112.822
R2378 w_570_7310.n127 w_570_7310.t14 112.822
R2379 w_570_7310.n127 w_570_7310.t25 112.822
R2380 w_570_7310.n308 w_570_7310.t29 112.822
R2381 w_570_7310.n308 w_570_7310.t10 112.822
R2382 w_570_7310.n203 w_570_7310.t12 112.822
R2383 w_570_7310.n366 w_570_7310.n363 20.092
R2384 w_570_7310.n424 w_570_7310.n423 16.607
R2385 w_570_7310.n276 w_570_7310.n275 16.289
R2386 w_570_7310.n126 w_570_7310.n125 16.289
R2387 w_570_7310.n51 w_570_7310.n50 16.289
R2388 w_570_7310.n500 w_570_7310.n499 16.288
R2389 w_570_7310.n211 w_570_7310.n207 12.923
R2390 w_570_7310.n429 w_570_7310.n425 12.641
R2391 w_570_7310.n8 w_570_7310.n4 12.629
R2392 w_570_7310.n60 w_570_7310.n56 12.629
R2393 w_570_7310.n135 w_570_7310.n131 12.629
R2394 w_570_7310.n281 w_570_7310.n277 12.629
R2395 w_570_7310.n201 w_570_7310.n200 12.369
R2396 w_570_7310.n431 w_570_7310.n430 9.3
R2397 w_570_7310.n437 w_570_7310.n436 9.3
R2398 w_570_7310.n443 w_570_7310.n442 9.3
R2399 w_570_7310.n449 w_570_7310.n448 9.3
R2400 w_570_7310.n455 w_570_7310.n454 9.3
R2401 w_570_7310.n467 w_570_7310.n466 9.3
R2402 w_570_7310.n473 w_570_7310.n472 9.3
R2403 w_570_7310.n479 w_570_7310.n478 9.3
R2404 w_570_7310.n485 w_570_7310.n484 9.3
R2405 w_570_7310.n491 w_570_7310.n490 9.3
R2406 w_570_7310.n496 w_570_7310.n495 9.3
R2407 w_570_7310.n62 w_570_7310.n61 9.3
R2408 w_570_7310.n68 w_570_7310.n67 9.3
R2409 w_570_7310.n74 w_570_7310.n73 9.3
R2410 w_570_7310.n80 w_570_7310.n79 9.3
R2411 w_570_7310.n86 w_570_7310.n85 9.3
R2412 w_570_7310.n94 w_570_7310.n93 9.3
R2413 w_570_7310.n100 w_570_7310.n99 9.3
R2414 w_570_7310.n106 w_570_7310.n105 9.3
R2415 w_570_7310.n112 w_570_7310.n111 9.3
R2416 w_570_7310.n118 w_570_7310.n117 9.3
R2417 w_570_7310.n123 w_570_7310.n122 9.3
R2418 w_570_7310.n137 w_570_7310.n136 9.3
R2419 w_570_7310.n143 w_570_7310.n142 9.3
R2420 w_570_7310.n149 w_570_7310.n148 9.3
R2421 w_570_7310.n155 w_570_7310.n154 9.3
R2422 w_570_7310.n161 w_570_7310.n160 9.3
R2423 w_570_7310.n169 w_570_7310.n168 9.3
R2424 w_570_7310.n175 w_570_7310.n174 9.3
R2425 w_570_7310.n181 w_570_7310.n180 9.3
R2426 w_570_7310.n187 w_570_7310.n186 9.3
R2427 w_570_7310.n193 w_570_7310.n192 9.3
R2428 w_570_7310.n198 w_570_7310.n197 9.3
R2429 w_570_7310.n273 w_570_7310.n272 9.3
R2430 w_570_7310.n213 w_570_7310.n212 9.3
R2431 w_570_7310.n219 w_570_7310.n218 9.3
R2432 w_570_7310.n225 w_570_7310.n224 9.3
R2433 w_570_7310.n231 w_570_7310.n230 9.3
R2434 w_570_7310.n237 w_570_7310.n236 9.3
R2435 w_570_7310.n245 w_570_7310.n244 9.3
R2436 w_570_7310.n251 w_570_7310.n250 9.3
R2437 w_570_7310.n257 w_570_7310.n256 9.3
R2438 w_570_7310.n263 w_570_7310.n262 9.3
R2439 w_570_7310.n268 w_570_7310.n267 9.3
R2440 w_570_7310.n283 w_570_7310.n282 9.3
R2441 w_570_7310.n289 w_570_7310.n288 9.3
R2442 w_570_7310.n295 w_570_7310.n294 9.3
R2443 w_570_7310.n301 w_570_7310.n300 9.3
R2444 w_570_7310.n307 w_570_7310.n306 9.3
R2445 w_570_7310.n319 w_570_7310.n318 9.3
R2446 w_570_7310.n325 w_570_7310.n324 9.3
R2447 w_570_7310.n331 w_570_7310.n330 9.3
R2448 w_570_7310.n337 w_570_7310.n336 9.3
R2449 w_570_7310.n343 w_570_7310.n342 9.3
R2450 w_570_7310.n348 w_570_7310.n347 9.3
R2451 w_570_7310.n287 w_570_7310.n286 9.3
R2452 w_570_7310.n293 w_570_7310.n292 9.3
R2453 w_570_7310.n299 w_570_7310.n298 9.3
R2454 w_570_7310.n305 w_570_7310.n304 9.3
R2455 w_570_7310.n323 w_570_7310.n322 9.3
R2456 w_570_7310.n329 w_570_7310.n328 9.3
R2457 w_570_7310.n335 w_570_7310.n334 9.3
R2458 w_570_7310.n341 w_570_7310.n340 9.3
R2459 w_570_7310.n346 w_570_7310.n345 9.3
R2460 w_570_7310.n141 w_570_7310.n140 9.3
R2461 w_570_7310.n147 w_570_7310.n146 9.3
R2462 w_570_7310.n153 w_570_7310.n152 9.3
R2463 w_570_7310.n159 w_570_7310.n158 9.3
R2464 w_570_7310.n173 w_570_7310.n172 9.3
R2465 w_570_7310.n179 w_570_7310.n178 9.3
R2466 w_570_7310.n185 w_570_7310.n184 9.3
R2467 w_570_7310.n191 w_570_7310.n190 9.3
R2468 w_570_7310.n196 w_570_7310.n195 9.3
R2469 w_570_7310.n66 w_570_7310.n65 9.3
R2470 w_570_7310.n72 w_570_7310.n71 9.3
R2471 w_570_7310.n78 w_570_7310.n77 9.3
R2472 w_570_7310.n84 w_570_7310.n83 9.3
R2473 w_570_7310.n98 w_570_7310.n97 9.3
R2474 w_570_7310.n104 w_570_7310.n103 9.3
R2475 w_570_7310.n110 w_570_7310.n109 9.3
R2476 w_570_7310.n116 w_570_7310.n115 9.3
R2477 w_570_7310.n121 w_570_7310.n120 9.3
R2478 w_570_7310.n435 w_570_7310.n434 9.3
R2479 w_570_7310.n441 w_570_7310.n440 9.3
R2480 w_570_7310.n447 w_570_7310.n446 9.3
R2481 w_570_7310.n453 w_570_7310.n452 9.3
R2482 w_570_7310.n471 w_570_7310.n470 9.3
R2483 w_570_7310.n477 w_570_7310.n476 9.3
R2484 w_570_7310.n483 w_570_7310.n482 9.3
R2485 w_570_7310.n489 w_570_7310.n488 9.3
R2486 w_570_7310.n494 w_570_7310.n493 9.3
R2487 w_570_7310.n217 w_570_7310.n216 9.3
R2488 w_570_7310.n223 w_570_7310.n222 9.3
R2489 w_570_7310.n229 w_570_7310.n228 9.3
R2490 w_570_7310.n235 w_570_7310.n234 9.3
R2491 w_570_7310.n249 w_570_7310.n248 9.3
R2492 w_570_7310.n255 w_570_7310.n254 9.3
R2493 w_570_7310.n261 w_570_7310.n260 9.3
R2494 w_570_7310.n266 w_570_7310.n265 9.3
R2495 w_570_7310.n271 w_570_7310.n270 9.3
R2496 w_570_7310.n368 w_570_7310.n367 9.3
R2497 w_570_7310.n371 w_570_7310.n370 9.3
R2498 w_570_7310.n373 w_570_7310.n372 9.3
R2499 w_570_7310.n376 w_570_7310.n375 9.3
R2500 w_570_7310.n378 w_570_7310.n377 9.3
R2501 w_570_7310.n381 w_570_7310.n380 9.3
R2502 w_570_7310.n383 w_570_7310.n382 9.3
R2503 w_570_7310.n386 w_570_7310.n385 9.3
R2504 w_570_7310.n388 w_570_7310.n387 9.3
R2505 w_570_7310.n395 w_570_7310.n394 9.3
R2506 w_570_7310.n398 w_570_7310.n397 9.3
R2507 w_570_7310.n400 w_570_7310.n399 9.3
R2508 w_570_7310.n403 w_570_7310.n402 9.3
R2509 w_570_7310.n405 w_570_7310.n404 9.3
R2510 w_570_7310.n408 w_570_7310.n407 9.3
R2511 w_570_7310.n410 w_570_7310.n409 9.3
R2512 w_570_7310.n413 w_570_7310.n412 9.3
R2513 w_570_7310.n415 w_570_7310.n414 9.3
R2514 w_570_7310.n418 w_570_7310.n417 9.3
R2515 w_570_7310.n420 w_570_7310.n419 9.3
R2516 w_570_7310.n10 w_570_7310.n9 9.3
R2517 w_570_7310.n14 w_570_7310.n13 9.3
R2518 w_570_7310.n16 w_570_7310.n15 9.3
R2519 w_570_7310.n20 w_570_7310.n19 9.3
R2520 w_570_7310.n22 w_570_7310.n21 9.3
R2521 w_570_7310.n26 w_570_7310.n25 9.3
R2522 w_570_7310.n28 w_570_7310.n27 9.3
R2523 w_570_7310.n32 w_570_7310.n31 9.3
R2524 w_570_7310.n34 w_570_7310.n33 9.3
R2525 w_570_7310.n532 w_570_7310.n531 9.3
R2526 w_570_7310.n530 w_570_7310.n529 9.3
R2527 w_570_7310.n526 w_570_7310.n525 9.3
R2528 w_570_7310.n524 w_570_7310.n523 9.3
R2529 w_570_7310.n520 w_570_7310.n519 9.3
R2530 w_570_7310.n518 w_570_7310.n517 9.3
R2531 w_570_7310.n514 w_570_7310.n513 9.3
R2532 w_570_7310.n512 w_570_7310.n511 9.3
R2533 w_570_7310.n508 w_570_7310.n507 9.3
R2534 w_570_7310.n506 w_570_7310.n505 9.3
R2535 w_570_7310.n503 w_570_7310.n502 9.3
R2536 w_570_7310.n280 w_570_7310.n279 8.855
R2537 w_570_7310.n286 w_570_7310.n285 8.855
R2538 w_570_7310.n292 w_570_7310.n291 8.855
R2539 w_570_7310.n298 w_570_7310.n297 8.855
R2540 w_570_7310.n304 w_570_7310.n303 8.855
R2541 w_570_7310.n311 w_570_7310.n310 8.855
R2542 w_570_7310.n316 w_570_7310.n315 8.855
R2543 w_570_7310.n322 w_570_7310.n321 8.855
R2544 w_570_7310.n328 w_570_7310.n327 8.855
R2545 w_570_7310.n334 w_570_7310.n333 8.855
R2546 w_570_7310.n340 w_570_7310.n339 8.855
R2547 w_570_7310.n345 w_570_7310.n344 8.855
R2548 w_570_7310.n134 w_570_7310.n133 8.855
R2549 w_570_7310.n140 w_570_7310.n139 8.855
R2550 w_570_7310.n146 w_570_7310.n145 8.855
R2551 w_570_7310.n152 w_570_7310.n151 8.855
R2552 w_570_7310.n158 w_570_7310.n157 8.855
R2553 w_570_7310.n130 w_570_7310.n129 8.855
R2554 w_570_7310.n166 w_570_7310.n165 8.855
R2555 w_570_7310.n172 w_570_7310.n171 8.855
R2556 w_570_7310.n178 w_570_7310.n177 8.855
R2557 w_570_7310.n184 w_570_7310.n183 8.855
R2558 w_570_7310.n190 w_570_7310.n189 8.855
R2559 w_570_7310.n195 w_570_7310.n194 8.855
R2560 w_570_7310.n59 w_570_7310.n58 8.855
R2561 w_570_7310.n65 w_570_7310.n64 8.855
R2562 w_570_7310.n71 w_570_7310.n70 8.855
R2563 w_570_7310.n77 w_570_7310.n76 8.855
R2564 w_570_7310.n83 w_570_7310.n82 8.855
R2565 w_570_7310.n55 w_570_7310.n54 8.855
R2566 w_570_7310.n91 w_570_7310.n90 8.855
R2567 w_570_7310.n97 w_570_7310.n96 8.855
R2568 w_570_7310.n103 w_570_7310.n102 8.855
R2569 w_570_7310.n109 w_570_7310.n108 8.855
R2570 w_570_7310.n115 w_570_7310.n114 8.855
R2571 w_570_7310.n120 w_570_7310.n119 8.855
R2572 w_570_7310.n7 w_570_7310.n6 8.855
R2573 w_570_7310.n428 w_570_7310.n427 8.855
R2574 w_570_7310.n434 w_570_7310.n433 8.855
R2575 w_570_7310.n440 w_570_7310.n439 8.855
R2576 w_570_7310.n446 w_570_7310.n445 8.855
R2577 w_570_7310.n452 w_570_7310.n451 8.855
R2578 w_570_7310.n459 w_570_7310.n458 8.855
R2579 w_570_7310.n464 w_570_7310.n463 8.855
R2580 w_570_7310.n470 w_570_7310.n469 8.855
R2581 w_570_7310.n476 w_570_7310.n475 8.855
R2582 w_570_7310.n482 w_570_7310.n481 8.855
R2583 w_570_7310.n488 w_570_7310.n487 8.855
R2584 w_570_7310.n493 w_570_7310.n492 8.855
R2585 w_570_7310.n210 w_570_7310.n209 8.855
R2586 w_570_7310.n216 w_570_7310.n215 8.855
R2587 w_570_7310.n222 w_570_7310.n221 8.855
R2588 w_570_7310.n228 w_570_7310.n227 8.855
R2589 w_570_7310.n234 w_570_7310.n233 8.855
R2590 w_570_7310.n240 w_570_7310.n239 8.855
R2591 w_570_7310.n206 w_570_7310.n205 8.855
R2592 w_570_7310.n248 w_570_7310.n247 8.855
R2593 w_570_7310.n254 w_570_7310.n253 8.855
R2594 w_570_7310.n260 w_570_7310.n259 8.855
R2595 w_570_7310.n265 w_570_7310.n264 8.855
R2596 w_570_7310.n270 w_570_7310.n269 8.855
R2597 w_570_7310.n365 w_570_7310.n364 8.855
R2598 w_570_7310.n370 w_570_7310.n369 8.855
R2599 w_570_7310.n375 w_570_7310.n374 8.855
R2600 w_570_7310.n380 w_570_7310.n379 8.855
R2601 w_570_7310.n385 w_570_7310.n384 8.855
R2602 w_570_7310.n362 w_570_7310.n361 8.855
R2603 w_570_7310.n392 w_570_7310.n391 8.855
R2604 w_570_7310.n397 w_570_7310.n396 8.855
R2605 w_570_7310.n402 w_570_7310.n401 8.855
R2606 w_570_7310.n407 w_570_7310.n406 8.855
R2607 w_570_7310.n412 w_570_7310.n411 8.855
R2608 w_570_7310.n417 w_570_7310.n416 8.855
R2609 w_570_7310.n13 w_570_7310.n12 8.855
R2610 w_570_7310.n19 w_570_7310.n18 8.855
R2611 w_570_7310.n25 w_570_7310.n24 8.855
R2612 w_570_7310.n31 w_570_7310.n30 8.855
R2613 w_570_7310.n3 w_570_7310.n2 8.855
R2614 w_570_7310.n38 w_570_7310.n37 8.855
R2615 w_570_7310.n529 w_570_7310.n528 8.855
R2616 w_570_7310.n523 w_570_7310.n522 8.855
R2617 w_570_7310.n517 w_570_7310.n516 8.855
R2618 w_570_7310.n511 w_570_7310.n510 8.855
R2619 w_570_7310.n505 w_570_7310.n504 8.855
R2620 w_570_7310.n361 w_570_7310.n360 7.463
R2621 w_570_7310.n349 w_570_7310.n276 6.209
R2622 w_570_7310.n199 w_570_7310.n126 6.209
R2623 w_570_7310.n124 w_570_7310.n51 6.209
R2624 w_570_7310.n421 w_570_7310.n353 6.209
R2625 w_570_7310.n501 w_570_7310.n500 6.209
R2626 w_570_7310.n497 w_570_7310.n424 6.208
R2627 w_570_7310.n309 w_570_7310.n308 5.95
R2628 w_570_7310.n128 w_570_7310.n127 5.95
R2629 w_570_7310.n53 w_570_7310.n52 5.95
R2630 w_570_7310.n1 w_570_7310.n0 5.95
R2631 w_570_7310.n317 w_570_7310.n316 5.876
R2632 w_570_7310.n167 w_570_7310.n166 5.876
R2633 w_570_7310.n92 w_570_7310.n91 5.876
R2634 w_570_7310.n393 w_570_7310.n392 5.876
R2635 w_570_7310.n533 w_570_7310.n38 5.876
R2636 w_570_7310.n241 w_570_7310.n240 5.873
R2637 w_570_7310.n465 w_570_7310.n464 5.873
R2638 w_570_7310.n534 w_570_7310.t24 5.713
R2639 w_570_7310.n390 w_570_7310.t7 5.713
R2640 w_570_7310.n461 w_570_7310.t32 5.713
R2641 w_570_7310.n313 w_570_7310.t30 5.713
R2642 w_570_7310.n313 w_570_7310.t11 5.713
R2643 w_570_7310.n88 w_570_7310.t28 5.713
R2644 w_570_7310.n88 w_570_7310.t9 5.713
R2645 w_570_7310.n163 w_570_7310.t15 5.713
R2646 w_570_7310.n163 w_570_7310.t26 5.713
R2647 w_570_7310.n242 w_570_7310.t13 5.713
R2648 w_570_7310.n390 w_570_7310.t34 5.713
R2649 w_570_7310.t17 w_570_7310.n534 5.713
R2650 w_570_7310.n274 w_570_7310.n201 5.637
R2651 w_570_7310.n60 w_570_7310.n59 5.614
R2652 w_570_7310.n135 w_570_7310.n134 5.614
R2653 w_570_7310.n281 w_570_7310.n280 5.614
R2654 w_570_7310.n366 w_570_7310.n365 5.614
R2655 w_570_7310.n8 w_570_7310.n7 5.614
R2656 w_570_7310.n429 w_570_7310.n428 5.611
R2657 w_570_7310.n211 w_570_7310.n210 5.571
R2658 w_570_7310.n457 w_570_7310.n456 5.347
R2659 w_570_7310.n204 w_570_7310.n203 5.347
R2660 w_570_7310.n39 w_570_7310.t21 4.491
R2661 w_570_7310.n39 w_570_7310.t20 4.386
R2662 w_570_7310.n40 w_570_7310.t4 4.386
R2663 w_570_7310.n41 w_570_7310.t2 4.386
R2664 w_570_7310.n42 w_570_7310.t5 4.386
R2665 w_570_7310.n43 w_570_7310.t0 4.386
R2666 w_570_7310.n44 w_570_7310.t18 4.386
R2667 w_570_7310.n45 w_570_7310.t19 4.386
R2668 w_570_7310.n46 w_570_7310.t35 4.386
R2669 w_570_7310.n47 w_570_7310.t22 4.386
R2670 w_570_7310.n48 w_570_7310.t3 4.386
R2671 w_570_7310.n49 w_570_7310.t1 4.386
R2672 w_570_7310.n312 w_570_7310.n311 4.27
R2673 w_570_7310.n162 w_570_7310.n130 4.27
R2674 w_570_7310.n87 w_570_7310.n55 4.27
R2675 w_570_7310.n389 w_570_7310.n362 4.27
R2676 w_570_7310.n35 w_570_7310.n3 4.27
R2677 w_570_7310.n460 w_570_7310.n459 4.269
R2678 w_570_7310.n243 w_570_7310.n206 4.269
R2679 w_570_7310.n259 w_570_7310.n258 3.685
R2680 w_570_7310.n253 w_570_7310.n252 3.685
R2681 w_570_7310.n247 w_570_7310.n246 3.685
R2682 w_570_7310.n205 w_570_7310.n204 3.685
R2683 w_570_7310.n239 w_570_7310.n238 3.685
R2684 w_570_7310.n233 w_570_7310.n232 3.685
R2685 w_570_7310.n227 w_570_7310.n226 3.685
R2686 w_570_7310.n221 w_570_7310.n220 3.685
R2687 w_570_7310.n215 w_570_7310.n214 3.685
R2688 w_570_7310.n487 w_570_7310.n486 3.685
R2689 w_570_7310.n481 w_570_7310.n480 3.685
R2690 w_570_7310.n475 w_570_7310.n474 3.685
R2691 w_570_7310.n469 w_570_7310.n468 3.685
R2692 w_570_7310.n463 w_570_7310.n462 3.685
R2693 w_570_7310.n458 w_570_7310.n457 3.685
R2694 w_570_7310.n451 w_570_7310.n450 3.685
R2695 w_570_7310.n445 w_570_7310.n444 3.685
R2696 w_570_7310.n439 w_570_7310.n438 3.685
R2697 w_570_7310.n433 w_570_7310.n432 3.685
R2698 w_570_7310.n209 w_570_7310.n208 3.514
R2699 w_570_7310.n427 w_570_7310.n426 3.514
R2700 w_570_7310.n510 w_570_7310.n509 3.052
R2701 w_570_7310.n516 w_570_7310.n515 3.052
R2702 w_570_7310.n522 w_570_7310.n521 3.052
R2703 w_570_7310.n528 w_570_7310.n527 3.052
R2704 w_570_7310.n37 w_570_7310.n36 3.052
R2705 w_570_7310.n2 w_570_7310.n1 3.052
R2706 w_570_7310.n30 w_570_7310.n29 3.052
R2707 w_570_7310.n24 w_570_7310.n23 3.052
R2708 w_570_7310.n18 w_570_7310.n17 3.052
R2709 w_570_7310.n12 w_570_7310.n11 3.052
R2710 w_570_7310.n114 w_570_7310.n113 3.052
R2711 w_570_7310.n108 w_570_7310.n107 3.052
R2712 w_570_7310.n102 w_570_7310.n101 3.052
R2713 w_570_7310.n96 w_570_7310.n95 3.052
R2714 w_570_7310.n90 w_570_7310.n89 3.052
R2715 w_570_7310.n54 w_570_7310.n53 3.052
R2716 w_570_7310.n82 w_570_7310.n81 3.052
R2717 w_570_7310.n76 w_570_7310.n75 3.052
R2718 w_570_7310.n70 w_570_7310.n69 3.052
R2719 w_570_7310.n64 w_570_7310.n63 3.052
R2720 w_570_7310.n189 w_570_7310.n188 3.052
R2721 w_570_7310.n183 w_570_7310.n182 3.052
R2722 w_570_7310.n177 w_570_7310.n176 3.052
R2723 w_570_7310.n171 w_570_7310.n170 3.052
R2724 w_570_7310.n165 w_570_7310.n164 3.052
R2725 w_570_7310.n129 w_570_7310.n128 3.052
R2726 w_570_7310.n157 w_570_7310.n156 3.052
R2727 w_570_7310.n151 w_570_7310.n150 3.052
R2728 w_570_7310.n145 w_570_7310.n144 3.052
R2729 w_570_7310.n139 w_570_7310.n138 3.052
R2730 w_570_7310.n339 w_570_7310.n338 3.052
R2731 w_570_7310.n333 w_570_7310.n332 3.052
R2732 w_570_7310.n327 w_570_7310.n326 3.052
R2733 w_570_7310.n321 w_570_7310.n320 3.052
R2734 w_570_7310.n315 w_570_7310.n314 3.052
R2735 w_570_7310.n310 w_570_7310.n309 3.052
R2736 w_570_7310.n303 w_570_7310.n302 3.052
R2737 w_570_7310.n297 w_570_7310.n296 3.052
R2738 w_570_7310.n291 w_570_7310.n290 3.052
R2739 w_570_7310.n285 w_570_7310.n284 3.052
R2740 w_570_7310.n6 w_570_7310.n5 2.91
R2741 w_570_7310.n58 w_570_7310.n57 2.91
R2742 w_570_7310.n133 w_570_7310.n132 2.91
R2743 w_570_7310.n279 w_570_7310.n278 2.91
R2744 w_570_7310.n352 w_570_7310.n49 2.351
R2745 w_570_7310.n350 w_570_7310.n274 0.768
R2746 w_570_7310.n498 w_570_7310.n497 0.75
R2747 w_570_7310.n213 w_570_7310.n211 0.713
R2748 w_570_7310.n359 w_570_7310.n358 0.697
R2749 w_570_7310.n359 w_570_7310.n357 0.697
R2750 w_570_7310.n360 w_570_7310.n359 0.697
R2751 w_570_7310.n359 w_570_7310.n356 0.697
R2752 w_570_7310.n359 w_570_7310.n355 0.697
R2753 w_570_7310.n359 w_570_7310.n354 0.697
R2754 w_570_7310.n431 w_570_7310.n429 0.668
R2755 w_570_7310.n368 w_570_7310.n366 0.652
R2756 w_570_7310.n10 w_570_7310.n8 0.652
R2757 w_570_7310.n62 w_570_7310.n60 0.652
R2758 w_570_7310.n137 w_570_7310.n135 0.652
R2759 w_570_7310.n283 w_570_7310.n281 0.652
R2760 w_570_7310.n203 w_570_7310.n202 0.592
R2761 w_570_7310.n422 w_570_7310.n352 0.57
R2762 w_570_7310.n352 w_570_7310.n351 0.57
R2763 w_570_7310.n351 w_570_7310.n350 0.57
R2764 w_570_7310.n498 w_570_7310.n422 0.57
R2765 w_570_7310.n352 w_570_7310.n124 0.208
R2766 w_570_7310.n351 w_570_7310.n199 0.208
R2767 w_570_7310.n350 w_570_7310.n349 0.208
R2768 w_570_7310.n422 w_570_7310.n421 0.208
R2769 w_570_7310.n501 w_570_7310.n498 0.208
R2770 w_570_7310.n41 w_570_7310.n40 0.106
R2771 w_570_7310.n43 w_570_7310.n42 0.106
R2772 w_570_7310.n45 w_570_7310.n44 0.106
R2773 w_570_7310.n47 w_570_7310.n46 0.106
R2774 w_570_7310.n49 w_570_7310.n48 0.106
R2775 w_570_7310.n40 w_570_7310.n39 0.083
R2776 w_570_7310.n42 w_570_7310.n41 0.083
R2777 w_570_7310.n44 w_570_7310.n43 0.083
R2778 w_570_7310.n46 w_570_7310.n45 0.083
R2779 w_570_7310.n48 w_570_7310.n47 0.083
R2780 w_570_7310.n467 w_570_7310.n465 0.047
R2781 w_570_7310.n241 w_570_7310.n237 0.046
R2782 w_570_7310.n274 w_570_7310.n273 0.045
R2783 w_570_7310.n460 w_570_7310.n455 0.043
R2784 w_570_7310.n245 w_570_7310.n243 0.042
R2785 w_570_7310.n497 w_570_7310.n496 0.04
R2786 w_570_7310.n496 w_570_7310.n494 0.032
R2787 w_570_7310.n494 w_570_7310.n491 0.032
R2788 w_570_7310.n491 w_570_7310.n489 0.032
R2789 w_570_7310.n489 w_570_7310.n485 0.032
R2790 w_570_7310.n485 w_570_7310.n483 0.032
R2791 w_570_7310.n483 w_570_7310.n479 0.032
R2792 w_570_7310.n479 w_570_7310.n477 0.032
R2793 w_570_7310.n477 w_570_7310.n473 0.032
R2794 w_570_7310.n473 w_570_7310.n471 0.032
R2795 w_570_7310.n471 w_570_7310.n467 0.032
R2796 w_570_7310.n455 w_570_7310.n453 0.032
R2797 w_570_7310.n453 w_570_7310.n449 0.032
R2798 w_570_7310.n449 w_570_7310.n447 0.032
R2799 w_570_7310.n447 w_570_7310.n443 0.032
R2800 w_570_7310.n443 w_570_7310.n441 0.032
R2801 w_570_7310.n441 w_570_7310.n437 0.032
R2802 w_570_7310.n437 w_570_7310.n435 0.032
R2803 w_570_7310.n435 w_570_7310.n431 0.032
R2804 w_570_7310.n94 w_570_7310.n92 0.031
R2805 w_570_7310.n169 w_570_7310.n167 0.031
R2806 w_570_7310.n319 w_570_7310.n317 0.031
R2807 w_570_7310.n395 w_570_7310.n393 0.031
R2808 w_570_7310.n533 w_570_7310.n532 0.031
R2809 w_570_7310.n273 w_570_7310.n271 0.031
R2810 w_570_7310.n271 w_570_7310.n268 0.031
R2811 w_570_7310.n268 w_570_7310.n266 0.031
R2812 w_570_7310.n266 w_570_7310.n263 0.031
R2813 w_570_7310.n263 w_570_7310.n261 0.031
R2814 w_570_7310.n261 w_570_7310.n257 0.031
R2815 w_570_7310.n257 w_570_7310.n255 0.031
R2816 w_570_7310.n255 w_570_7310.n251 0.031
R2817 w_570_7310.n251 w_570_7310.n249 0.031
R2818 w_570_7310.n249 w_570_7310.n245 0.031
R2819 w_570_7310.n237 w_570_7310.n235 0.031
R2820 w_570_7310.n235 w_570_7310.n231 0.031
R2821 w_570_7310.n231 w_570_7310.n229 0.031
R2822 w_570_7310.n229 w_570_7310.n225 0.031
R2823 w_570_7310.n225 w_570_7310.n223 0.031
R2824 w_570_7310.n223 w_570_7310.n219 0.031
R2825 w_570_7310.n219 w_570_7310.n217 0.031
R2826 w_570_7310.n217 w_570_7310.n213 0.031
R2827 w_570_7310.n465 w_570_7310.n461 0.031
R2828 w_570_7310.n242 w_570_7310.n241 0.03
R2829 w_570_7310.n87 w_570_7310.n86 0.029
R2830 w_570_7310.n162 w_570_7310.n161 0.029
R2831 w_570_7310.n312 w_570_7310.n307 0.029
R2832 w_570_7310.n389 w_570_7310.n388 0.029
R2833 w_570_7310.n35 w_570_7310.n34 0.029
R2834 w_570_7310.n124 w_570_7310.n123 0.027
R2835 w_570_7310.n199 w_570_7310.n198 0.027
R2836 w_570_7310.n349 w_570_7310.n348 0.027
R2837 w_570_7310.n421 w_570_7310.n420 0.027
R2838 w_570_7310.n503 w_570_7310.n501 0.027
R2839 w_570_7310.n123 w_570_7310.n121 0.021
R2840 w_570_7310.n121 w_570_7310.n118 0.021
R2841 w_570_7310.n118 w_570_7310.n116 0.021
R2842 w_570_7310.n116 w_570_7310.n112 0.021
R2843 w_570_7310.n112 w_570_7310.n110 0.021
R2844 w_570_7310.n110 w_570_7310.n106 0.021
R2845 w_570_7310.n106 w_570_7310.n104 0.021
R2846 w_570_7310.n104 w_570_7310.n100 0.021
R2847 w_570_7310.n100 w_570_7310.n98 0.021
R2848 w_570_7310.n98 w_570_7310.n94 0.021
R2849 w_570_7310.n86 w_570_7310.n84 0.021
R2850 w_570_7310.n84 w_570_7310.n80 0.021
R2851 w_570_7310.n80 w_570_7310.n78 0.021
R2852 w_570_7310.n78 w_570_7310.n74 0.021
R2853 w_570_7310.n74 w_570_7310.n72 0.021
R2854 w_570_7310.n72 w_570_7310.n68 0.021
R2855 w_570_7310.n68 w_570_7310.n66 0.021
R2856 w_570_7310.n66 w_570_7310.n62 0.021
R2857 w_570_7310.n198 w_570_7310.n196 0.021
R2858 w_570_7310.n196 w_570_7310.n193 0.021
R2859 w_570_7310.n193 w_570_7310.n191 0.021
R2860 w_570_7310.n191 w_570_7310.n187 0.021
R2861 w_570_7310.n187 w_570_7310.n185 0.021
R2862 w_570_7310.n185 w_570_7310.n181 0.021
R2863 w_570_7310.n181 w_570_7310.n179 0.021
R2864 w_570_7310.n179 w_570_7310.n175 0.021
R2865 w_570_7310.n175 w_570_7310.n173 0.021
R2866 w_570_7310.n173 w_570_7310.n169 0.021
R2867 w_570_7310.n161 w_570_7310.n159 0.021
R2868 w_570_7310.n159 w_570_7310.n155 0.021
R2869 w_570_7310.n155 w_570_7310.n153 0.021
R2870 w_570_7310.n153 w_570_7310.n149 0.021
R2871 w_570_7310.n149 w_570_7310.n147 0.021
R2872 w_570_7310.n147 w_570_7310.n143 0.021
R2873 w_570_7310.n143 w_570_7310.n141 0.021
R2874 w_570_7310.n141 w_570_7310.n137 0.021
R2875 w_570_7310.n348 w_570_7310.n346 0.021
R2876 w_570_7310.n346 w_570_7310.n343 0.021
R2877 w_570_7310.n343 w_570_7310.n341 0.021
R2878 w_570_7310.n341 w_570_7310.n337 0.021
R2879 w_570_7310.n337 w_570_7310.n335 0.021
R2880 w_570_7310.n335 w_570_7310.n331 0.021
R2881 w_570_7310.n331 w_570_7310.n329 0.021
R2882 w_570_7310.n329 w_570_7310.n325 0.021
R2883 w_570_7310.n325 w_570_7310.n323 0.021
R2884 w_570_7310.n323 w_570_7310.n319 0.021
R2885 w_570_7310.n307 w_570_7310.n305 0.021
R2886 w_570_7310.n305 w_570_7310.n301 0.021
R2887 w_570_7310.n301 w_570_7310.n299 0.021
R2888 w_570_7310.n299 w_570_7310.n295 0.021
R2889 w_570_7310.n295 w_570_7310.n293 0.021
R2890 w_570_7310.n293 w_570_7310.n289 0.021
R2891 w_570_7310.n289 w_570_7310.n287 0.021
R2892 w_570_7310.n287 w_570_7310.n283 0.021
R2893 w_570_7310.n420 w_570_7310.n418 0.021
R2894 w_570_7310.n418 w_570_7310.n415 0.021
R2895 w_570_7310.n415 w_570_7310.n413 0.021
R2896 w_570_7310.n413 w_570_7310.n410 0.021
R2897 w_570_7310.n410 w_570_7310.n408 0.021
R2898 w_570_7310.n408 w_570_7310.n405 0.021
R2899 w_570_7310.n405 w_570_7310.n403 0.021
R2900 w_570_7310.n403 w_570_7310.n400 0.021
R2901 w_570_7310.n400 w_570_7310.n398 0.021
R2902 w_570_7310.n398 w_570_7310.n395 0.021
R2903 w_570_7310.n388 w_570_7310.n386 0.021
R2904 w_570_7310.n386 w_570_7310.n383 0.021
R2905 w_570_7310.n383 w_570_7310.n381 0.021
R2906 w_570_7310.n381 w_570_7310.n378 0.021
R2907 w_570_7310.n378 w_570_7310.n376 0.021
R2908 w_570_7310.n376 w_570_7310.n373 0.021
R2909 w_570_7310.n373 w_570_7310.n371 0.021
R2910 w_570_7310.n371 w_570_7310.n368 0.021
R2911 w_570_7310.n506 w_570_7310.n503 0.021
R2912 w_570_7310.n508 w_570_7310.n506 0.021
R2913 w_570_7310.n512 w_570_7310.n508 0.021
R2914 w_570_7310.n514 w_570_7310.n512 0.021
R2915 w_570_7310.n518 w_570_7310.n514 0.021
R2916 w_570_7310.n520 w_570_7310.n518 0.021
R2917 w_570_7310.n524 w_570_7310.n520 0.021
R2918 w_570_7310.n526 w_570_7310.n524 0.021
R2919 w_570_7310.n530 w_570_7310.n526 0.021
R2920 w_570_7310.n532 w_570_7310.n530 0.021
R2921 w_570_7310.n34 w_570_7310.n32 0.021
R2922 w_570_7310.n32 w_570_7310.n28 0.021
R2923 w_570_7310.n28 w_570_7310.n26 0.021
R2924 w_570_7310.n26 w_570_7310.n22 0.021
R2925 w_570_7310.n22 w_570_7310.n20 0.021
R2926 w_570_7310.n20 w_570_7310.n16 0.021
R2927 w_570_7310.n16 w_570_7310.n14 0.021
R2928 w_570_7310.n14 w_570_7310.n10 0.021
R2929 w_570_7310.n534 w_570_7310.n533 0.021
R2930 w_570_7310.n92 w_570_7310.n88 0.021
R2931 w_570_7310.n167 w_570_7310.n163 0.021
R2932 w_570_7310.n317 w_570_7310.n313 0.021
R2933 w_570_7310.n393 w_570_7310.n390 0.021
R2934 w_570_7310.n461 w_570_7310.n460 0.009
R2935 w_570_7310.n243 w_570_7310.n242 0.009
R2936 w_570_7310.n534 w_570_7310.n35 0.006
R2937 w_570_7310.n88 w_570_7310.n87 0.006
R2938 w_570_7310.n163 w_570_7310.n162 0.006
R2939 w_570_7310.n313 w_570_7310.n312 0.006
R2940 w_570_7310.n390 w_570_7310.n389 0.006
R2941 w_6940_7310.n329 w_6940_7310.t28 112.822
R2942 w_6940_7310.n373 w_6940_7310.t4 112.822
R2943 w_6940_7310.n373 w_6940_7310.t2 112.822
R2944 w_6940_7310.n480 w_6940_7310.t22 112.822
R2945 w_6940_7310.n480 w_6940_7310.t12 112.822
R2946 w_6940_7310.n6 w_6940_7310.t26 112.822
R2947 w_6940_7310.n6 w_6940_7310.t10 112.822
R2948 w_6940_7310.n71 w_6940_7310.t24 112.822
R2949 w_6940_7310.n71 w_6940_7310.t8 112.822
R2950 w_6940_7310.n252 w_6940_7310.t6 112.822
R2951 w_6940_7310.n252 w_6940_7310.t0 112.822
R2952 w_6940_7310.n147 w_6940_7310.t20 112.822
R2953 w_6940_7310.n13 w_6940_7310.n10 20.092
R2954 w_6940_7310.n297 w_6940_7310.n296 16.607
R2955 w_6940_7310.n220 w_6940_7310.n219 16.289
R2956 w_6940_7310.n70 w_6940_7310.n69 16.289
R2957 w_6940_7310.n448 w_6940_7310.n447 16.289
R2958 w_6940_7310.n372 w_6940_7310.n371 16.289
R2959 w_6940_7310.n155 w_6940_7310.n151 12.923
R2960 w_6940_7310.n302 w_6940_7310.n298 12.641
R2961 w_6940_7310.n381 w_6940_7310.n377 12.629
R2962 w_6940_7310.n453 w_6940_7310.n449 12.629
R2963 w_6940_7310.n79 w_6940_7310.n75 12.629
R2964 w_6940_7310.n225 w_6940_7310.n221 12.629
R2965 w_6940_7310.n145 w_6940_7310.n144 12.369
R2966 w_6940_7310.n304 w_6940_7310.n303 9.3
R2967 w_6940_7310.n310 w_6940_7310.n309 9.3
R2968 w_6940_7310.n316 w_6940_7310.n315 9.3
R2969 w_6940_7310.n322 w_6940_7310.n321 9.3
R2970 w_6940_7310.n328 w_6940_7310.n327 9.3
R2971 w_6940_7310.n340 w_6940_7310.n339 9.3
R2972 w_6940_7310.n346 w_6940_7310.n345 9.3
R2973 w_6940_7310.n352 w_6940_7310.n351 9.3
R2974 w_6940_7310.n358 w_6940_7310.n357 9.3
R2975 w_6940_7310.n364 w_6940_7310.n363 9.3
R2976 w_6940_7310.n369 w_6940_7310.n368 9.3
R2977 w_6940_7310.n383 w_6940_7310.n382 9.3
R2978 w_6940_7310.n389 w_6940_7310.n388 9.3
R2979 w_6940_7310.n395 w_6940_7310.n394 9.3
R2980 w_6940_7310.n401 w_6940_7310.n400 9.3
R2981 w_6940_7310.n407 w_6940_7310.n406 9.3
R2982 w_6940_7310.n415 w_6940_7310.n414 9.3
R2983 w_6940_7310.n421 w_6940_7310.n420 9.3
R2984 w_6940_7310.n427 w_6940_7310.n426 9.3
R2985 w_6940_7310.n433 w_6940_7310.n432 9.3
R2986 w_6940_7310.n439 w_6940_7310.n438 9.3
R2987 w_6940_7310.n444 w_6940_7310.n443 9.3
R2988 w_6940_7310.n455 w_6940_7310.n454 9.3
R2989 w_6940_7310.n461 w_6940_7310.n460 9.3
R2990 w_6940_7310.n467 w_6940_7310.n466 9.3
R2991 w_6940_7310.n473 w_6940_7310.n472 9.3
R2992 w_6940_7310.n479 w_6940_7310.n478 9.3
R2993 w_6940_7310.n491 w_6940_7310.n490 9.3
R2994 w_6940_7310.n497 w_6940_7310.n496 9.3
R2995 w_6940_7310.n503 w_6940_7310.n502 9.3
R2996 w_6940_7310.n509 w_6940_7310.n508 9.3
R2997 w_6940_7310.n515 w_6940_7310.n514 9.3
R2998 w_6940_7310.n520 w_6940_7310.n519 9.3
R2999 w_6940_7310.n81 w_6940_7310.n80 9.3
R3000 w_6940_7310.n87 w_6940_7310.n86 9.3
R3001 w_6940_7310.n93 w_6940_7310.n92 9.3
R3002 w_6940_7310.n99 w_6940_7310.n98 9.3
R3003 w_6940_7310.n105 w_6940_7310.n104 9.3
R3004 w_6940_7310.n113 w_6940_7310.n112 9.3
R3005 w_6940_7310.n119 w_6940_7310.n118 9.3
R3006 w_6940_7310.n125 w_6940_7310.n124 9.3
R3007 w_6940_7310.n131 w_6940_7310.n130 9.3
R3008 w_6940_7310.n137 w_6940_7310.n136 9.3
R3009 w_6940_7310.n142 w_6940_7310.n141 9.3
R3010 w_6940_7310.n217 w_6940_7310.n216 9.3
R3011 w_6940_7310.n157 w_6940_7310.n156 9.3
R3012 w_6940_7310.n163 w_6940_7310.n162 9.3
R3013 w_6940_7310.n169 w_6940_7310.n168 9.3
R3014 w_6940_7310.n175 w_6940_7310.n174 9.3
R3015 w_6940_7310.n181 w_6940_7310.n180 9.3
R3016 w_6940_7310.n189 w_6940_7310.n188 9.3
R3017 w_6940_7310.n195 w_6940_7310.n194 9.3
R3018 w_6940_7310.n201 w_6940_7310.n200 9.3
R3019 w_6940_7310.n207 w_6940_7310.n206 9.3
R3020 w_6940_7310.n212 w_6940_7310.n211 9.3
R3021 w_6940_7310.n227 w_6940_7310.n226 9.3
R3022 w_6940_7310.n233 w_6940_7310.n232 9.3
R3023 w_6940_7310.n239 w_6940_7310.n238 9.3
R3024 w_6940_7310.n245 w_6940_7310.n244 9.3
R3025 w_6940_7310.n251 w_6940_7310.n250 9.3
R3026 w_6940_7310.n263 w_6940_7310.n262 9.3
R3027 w_6940_7310.n269 w_6940_7310.n268 9.3
R3028 w_6940_7310.n275 w_6940_7310.n274 9.3
R3029 w_6940_7310.n281 w_6940_7310.n280 9.3
R3030 w_6940_7310.n287 w_6940_7310.n286 9.3
R3031 w_6940_7310.n292 w_6940_7310.n291 9.3
R3032 w_6940_7310.n231 w_6940_7310.n230 9.3
R3033 w_6940_7310.n237 w_6940_7310.n236 9.3
R3034 w_6940_7310.n243 w_6940_7310.n242 9.3
R3035 w_6940_7310.n249 w_6940_7310.n248 9.3
R3036 w_6940_7310.n267 w_6940_7310.n266 9.3
R3037 w_6940_7310.n273 w_6940_7310.n272 9.3
R3038 w_6940_7310.n279 w_6940_7310.n278 9.3
R3039 w_6940_7310.n285 w_6940_7310.n284 9.3
R3040 w_6940_7310.n290 w_6940_7310.n289 9.3
R3041 w_6940_7310.n85 w_6940_7310.n84 9.3
R3042 w_6940_7310.n91 w_6940_7310.n90 9.3
R3043 w_6940_7310.n97 w_6940_7310.n96 9.3
R3044 w_6940_7310.n103 w_6940_7310.n102 9.3
R3045 w_6940_7310.n117 w_6940_7310.n116 9.3
R3046 w_6940_7310.n123 w_6940_7310.n122 9.3
R3047 w_6940_7310.n129 w_6940_7310.n128 9.3
R3048 w_6940_7310.n135 w_6940_7310.n134 9.3
R3049 w_6940_7310.n140 w_6940_7310.n139 9.3
R3050 w_6940_7310.n459 w_6940_7310.n458 9.3
R3051 w_6940_7310.n465 w_6940_7310.n464 9.3
R3052 w_6940_7310.n471 w_6940_7310.n470 9.3
R3053 w_6940_7310.n477 w_6940_7310.n476 9.3
R3054 w_6940_7310.n495 w_6940_7310.n494 9.3
R3055 w_6940_7310.n501 w_6940_7310.n500 9.3
R3056 w_6940_7310.n507 w_6940_7310.n506 9.3
R3057 w_6940_7310.n513 w_6940_7310.n512 9.3
R3058 w_6940_7310.n518 w_6940_7310.n517 9.3
R3059 w_6940_7310.n387 w_6940_7310.n386 9.3
R3060 w_6940_7310.n393 w_6940_7310.n392 9.3
R3061 w_6940_7310.n399 w_6940_7310.n398 9.3
R3062 w_6940_7310.n405 w_6940_7310.n404 9.3
R3063 w_6940_7310.n419 w_6940_7310.n418 9.3
R3064 w_6940_7310.n425 w_6940_7310.n424 9.3
R3065 w_6940_7310.n431 w_6940_7310.n430 9.3
R3066 w_6940_7310.n437 w_6940_7310.n436 9.3
R3067 w_6940_7310.n442 w_6940_7310.n441 9.3
R3068 w_6940_7310.n308 w_6940_7310.n307 9.3
R3069 w_6940_7310.n314 w_6940_7310.n313 9.3
R3070 w_6940_7310.n320 w_6940_7310.n319 9.3
R3071 w_6940_7310.n326 w_6940_7310.n325 9.3
R3072 w_6940_7310.n344 w_6940_7310.n343 9.3
R3073 w_6940_7310.n350 w_6940_7310.n349 9.3
R3074 w_6940_7310.n356 w_6940_7310.n355 9.3
R3075 w_6940_7310.n362 w_6940_7310.n361 9.3
R3076 w_6940_7310.n367 w_6940_7310.n366 9.3
R3077 w_6940_7310.n161 w_6940_7310.n160 9.3
R3078 w_6940_7310.n167 w_6940_7310.n166 9.3
R3079 w_6940_7310.n173 w_6940_7310.n172 9.3
R3080 w_6940_7310.n179 w_6940_7310.n178 9.3
R3081 w_6940_7310.n193 w_6940_7310.n192 9.3
R3082 w_6940_7310.n199 w_6940_7310.n198 9.3
R3083 w_6940_7310.n205 w_6940_7310.n204 9.3
R3084 w_6940_7310.n210 w_6940_7310.n209 9.3
R3085 w_6940_7310.n215 w_6940_7310.n214 9.3
R3086 w_6940_7310.n15 w_6940_7310.n14 9.3
R3087 w_6940_7310.n18 w_6940_7310.n17 9.3
R3088 w_6940_7310.n20 w_6940_7310.n19 9.3
R3089 w_6940_7310.n23 w_6940_7310.n22 9.3
R3090 w_6940_7310.n25 w_6940_7310.n24 9.3
R3091 w_6940_7310.n28 w_6940_7310.n27 9.3
R3092 w_6940_7310.n30 w_6940_7310.n29 9.3
R3093 w_6940_7310.n33 w_6940_7310.n32 9.3
R3094 w_6940_7310.n35 w_6940_7310.n34 9.3
R3095 w_6940_7310.n42 w_6940_7310.n41 9.3
R3096 w_6940_7310.n45 w_6940_7310.n44 9.3
R3097 w_6940_7310.n47 w_6940_7310.n46 9.3
R3098 w_6940_7310.n50 w_6940_7310.n49 9.3
R3099 w_6940_7310.n52 w_6940_7310.n51 9.3
R3100 w_6940_7310.n55 w_6940_7310.n54 9.3
R3101 w_6940_7310.n57 w_6940_7310.n56 9.3
R3102 w_6940_7310.n60 w_6940_7310.n59 9.3
R3103 w_6940_7310.n62 w_6940_7310.n61 9.3
R3104 w_6940_7310.n65 w_6940_7310.n64 9.3
R3105 w_6940_7310.n67 w_6940_7310.n66 9.3
R3106 w_6940_7310.n224 w_6940_7310.n223 8.855
R3107 w_6940_7310.n230 w_6940_7310.n229 8.855
R3108 w_6940_7310.n236 w_6940_7310.n235 8.855
R3109 w_6940_7310.n242 w_6940_7310.n241 8.855
R3110 w_6940_7310.n248 w_6940_7310.n247 8.855
R3111 w_6940_7310.n255 w_6940_7310.n254 8.855
R3112 w_6940_7310.n260 w_6940_7310.n259 8.855
R3113 w_6940_7310.n266 w_6940_7310.n265 8.855
R3114 w_6940_7310.n272 w_6940_7310.n271 8.855
R3115 w_6940_7310.n278 w_6940_7310.n277 8.855
R3116 w_6940_7310.n284 w_6940_7310.n283 8.855
R3117 w_6940_7310.n289 w_6940_7310.n288 8.855
R3118 w_6940_7310.n78 w_6940_7310.n77 8.855
R3119 w_6940_7310.n84 w_6940_7310.n83 8.855
R3120 w_6940_7310.n90 w_6940_7310.n89 8.855
R3121 w_6940_7310.n96 w_6940_7310.n95 8.855
R3122 w_6940_7310.n102 w_6940_7310.n101 8.855
R3123 w_6940_7310.n74 w_6940_7310.n73 8.855
R3124 w_6940_7310.n110 w_6940_7310.n109 8.855
R3125 w_6940_7310.n116 w_6940_7310.n115 8.855
R3126 w_6940_7310.n122 w_6940_7310.n121 8.855
R3127 w_6940_7310.n128 w_6940_7310.n127 8.855
R3128 w_6940_7310.n134 w_6940_7310.n133 8.855
R3129 w_6940_7310.n139 w_6940_7310.n138 8.855
R3130 w_6940_7310.n452 w_6940_7310.n451 8.855
R3131 w_6940_7310.n458 w_6940_7310.n457 8.855
R3132 w_6940_7310.n464 w_6940_7310.n463 8.855
R3133 w_6940_7310.n470 w_6940_7310.n469 8.855
R3134 w_6940_7310.n476 w_6940_7310.n475 8.855
R3135 w_6940_7310.n483 w_6940_7310.n482 8.855
R3136 w_6940_7310.n488 w_6940_7310.n487 8.855
R3137 w_6940_7310.n494 w_6940_7310.n493 8.855
R3138 w_6940_7310.n500 w_6940_7310.n499 8.855
R3139 w_6940_7310.n506 w_6940_7310.n505 8.855
R3140 w_6940_7310.n512 w_6940_7310.n511 8.855
R3141 w_6940_7310.n517 w_6940_7310.n516 8.855
R3142 w_6940_7310.n380 w_6940_7310.n379 8.855
R3143 w_6940_7310.n386 w_6940_7310.n385 8.855
R3144 w_6940_7310.n392 w_6940_7310.n391 8.855
R3145 w_6940_7310.n398 w_6940_7310.n397 8.855
R3146 w_6940_7310.n404 w_6940_7310.n403 8.855
R3147 w_6940_7310.n376 w_6940_7310.n375 8.855
R3148 w_6940_7310.n412 w_6940_7310.n411 8.855
R3149 w_6940_7310.n418 w_6940_7310.n417 8.855
R3150 w_6940_7310.n424 w_6940_7310.n423 8.855
R3151 w_6940_7310.n430 w_6940_7310.n429 8.855
R3152 w_6940_7310.n436 w_6940_7310.n435 8.855
R3153 w_6940_7310.n441 w_6940_7310.n440 8.855
R3154 w_6940_7310.n301 w_6940_7310.n300 8.855
R3155 w_6940_7310.n307 w_6940_7310.n306 8.855
R3156 w_6940_7310.n313 w_6940_7310.n312 8.855
R3157 w_6940_7310.n319 w_6940_7310.n318 8.855
R3158 w_6940_7310.n325 w_6940_7310.n324 8.855
R3159 w_6940_7310.n332 w_6940_7310.n331 8.855
R3160 w_6940_7310.n337 w_6940_7310.n336 8.855
R3161 w_6940_7310.n343 w_6940_7310.n342 8.855
R3162 w_6940_7310.n349 w_6940_7310.n348 8.855
R3163 w_6940_7310.n355 w_6940_7310.n354 8.855
R3164 w_6940_7310.n361 w_6940_7310.n360 8.855
R3165 w_6940_7310.n366 w_6940_7310.n365 8.855
R3166 w_6940_7310.n154 w_6940_7310.n153 8.855
R3167 w_6940_7310.n160 w_6940_7310.n159 8.855
R3168 w_6940_7310.n166 w_6940_7310.n165 8.855
R3169 w_6940_7310.n172 w_6940_7310.n171 8.855
R3170 w_6940_7310.n178 w_6940_7310.n177 8.855
R3171 w_6940_7310.n184 w_6940_7310.n183 8.855
R3172 w_6940_7310.n150 w_6940_7310.n149 8.855
R3173 w_6940_7310.n192 w_6940_7310.n191 8.855
R3174 w_6940_7310.n198 w_6940_7310.n197 8.855
R3175 w_6940_7310.n204 w_6940_7310.n203 8.855
R3176 w_6940_7310.n209 w_6940_7310.n208 8.855
R3177 w_6940_7310.n214 w_6940_7310.n213 8.855
R3178 w_6940_7310.n12 w_6940_7310.n11 8.855
R3179 w_6940_7310.n17 w_6940_7310.n16 8.855
R3180 w_6940_7310.n22 w_6940_7310.n21 8.855
R3181 w_6940_7310.n27 w_6940_7310.n26 8.855
R3182 w_6940_7310.n32 w_6940_7310.n31 8.855
R3183 w_6940_7310.n9 w_6940_7310.n8 8.855
R3184 w_6940_7310.n39 w_6940_7310.n38 8.855
R3185 w_6940_7310.n44 w_6940_7310.n43 8.855
R3186 w_6940_7310.n49 w_6940_7310.n48 8.855
R3187 w_6940_7310.n54 w_6940_7310.n53 8.855
R3188 w_6940_7310.n59 w_6940_7310.n58 8.855
R3189 w_6940_7310.n64 w_6940_7310.n63 8.855
R3190 w_6940_7310.n8 w_6940_7310.n7 7.463
R3191 w_6940_7310.n293 w_6940_7310.n220 6.209
R3192 w_6940_7310.n143 w_6940_7310.n70 6.209
R3193 w_6940_7310.n521 w_6940_7310.n448 6.209
R3194 w_6940_7310.n445 w_6940_7310.n372 6.209
R3195 w_6940_7310.n68 w_6940_7310.n0 6.209
R3196 w_6940_7310.n370 w_6940_7310.n297 6.208
R3197 w_6940_7310.n253 w_6940_7310.n252 5.95
R3198 w_6940_7310.n72 w_6940_7310.n71 5.95
R3199 w_6940_7310.n481 w_6940_7310.n480 5.95
R3200 w_6940_7310.n374 w_6940_7310.n373 5.95
R3201 w_6940_7310.n261 w_6940_7310.n260 5.876
R3202 w_6940_7310.n111 w_6940_7310.n110 5.876
R3203 w_6940_7310.n489 w_6940_7310.n488 5.876
R3204 w_6940_7310.n413 w_6940_7310.n412 5.876
R3205 w_6940_7310.n40 w_6940_7310.n39 5.876
R3206 w_6940_7310.n185 w_6940_7310.n184 5.873
R3207 w_6940_7310.n338 w_6940_7310.n337 5.873
R3208 w_6940_7310.n37 w_6940_7310.t27 5.713
R3209 w_6940_7310.n485 w_6940_7310.t23 5.713
R3210 w_6940_7310.n485 w_6940_7310.t13 5.713
R3211 w_6940_7310.n334 w_6940_7310.t29 5.713
R3212 w_6940_7310.n409 w_6940_7310.t5 5.713
R3213 w_6940_7310.n409 w_6940_7310.t3 5.713
R3214 w_6940_7310.n257 w_6940_7310.t7 5.713
R3215 w_6940_7310.n257 w_6940_7310.t1 5.713
R3216 w_6940_7310.n107 w_6940_7310.t25 5.713
R3217 w_6940_7310.n107 w_6940_7310.t9 5.713
R3218 w_6940_7310.n186 w_6940_7310.t21 5.713
R3219 w_6940_7310.n37 w_6940_7310.t11 5.713
R3220 w_6940_7310.n218 w_6940_7310.n145 5.637
R3221 w_6940_7310.n381 w_6940_7310.n380 5.614
R3222 w_6940_7310.n79 w_6940_7310.n78 5.614
R3223 w_6940_7310.n225 w_6940_7310.n224 5.614
R3224 w_6940_7310.n453 w_6940_7310.n452 5.614
R3225 w_6940_7310.n13 w_6940_7310.n12 5.614
R3226 w_6940_7310.n302 w_6940_7310.n301 5.611
R3227 w_6940_7310.n155 w_6940_7310.n154 5.571
R3228 w_6940_7310.n330 w_6940_7310.n329 5.347
R3229 w_6940_7310.n148 w_6940_7310.n147 5.347
R3230 w_6940_7310.n529 w_6940_7310.t32 4.491
R3231 w_6940_7310.n529 w_6940_7310.t34 4.386
R3232 w_6940_7310.n530 w_6940_7310.t18 4.386
R3233 w_6940_7310.n531 w_6940_7310.t14 4.386
R3234 w_6940_7310.n532 w_6940_7310.t33 4.386
R3235 w_6940_7310.n533 w_6940_7310.t35 4.386
R3236 w_6940_7310.n528 w_6940_7310.t16 4.386
R3237 w_6940_7310.n527 w_6940_7310.t30 4.386
R3238 w_6940_7310.n526 w_6940_7310.t31 4.386
R3239 w_6940_7310.n525 w_6940_7310.t15 4.386
R3240 w_6940_7310.n524 w_6940_7310.t17 4.386
R3241 w_6940_7310.t19 w_6940_7310.n534 4.385
R3242 w_6940_7310.n484 w_6940_7310.n483 4.27
R3243 w_6940_7310.n256 w_6940_7310.n255 4.27
R3244 w_6940_7310.n106 w_6940_7310.n74 4.27
R3245 w_6940_7310.n408 w_6940_7310.n376 4.27
R3246 w_6940_7310.n36 w_6940_7310.n9 4.27
R3247 w_6940_7310.n333 w_6940_7310.n332 4.269
R3248 w_6940_7310.n187 w_6940_7310.n150 4.269
R3249 w_6940_7310.n203 w_6940_7310.n202 3.685
R3250 w_6940_7310.n197 w_6940_7310.n196 3.685
R3251 w_6940_7310.n191 w_6940_7310.n190 3.685
R3252 w_6940_7310.n149 w_6940_7310.n148 3.685
R3253 w_6940_7310.n183 w_6940_7310.n182 3.685
R3254 w_6940_7310.n177 w_6940_7310.n176 3.685
R3255 w_6940_7310.n171 w_6940_7310.n170 3.685
R3256 w_6940_7310.n165 w_6940_7310.n164 3.685
R3257 w_6940_7310.n159 w_6940_7310.n158 3.685
R3258 w_6940_7310.n360 w_6940_7310.n359 3.685
R3259 w_6940_7310.n354 w_6940_7310.n353 3.685
R3260 w_6940_7310.n348 w_6940_7310.n347 3.685
R3261 w_6940_7310.n342 w_6940_7310.n341 3.685
R3262 w_6940_7310.n336 w_6940_7310.n335 3.685
R3263 w_6940_7310.n331 w_6940_7310.n330 3.685
R3264 w_6940_7310.n324 w_6940_7310.n323 3.685
R3265 w_6940_7310.n318 w_6940_7310.n317 3.685
R3266 w_6940_7310.n312 w_6940_7310.n311 3.685
R3267 w_6940_7310.n306 w_6940_7310.n305 3.685
R3268 w_6940_7310.n153 w_6940_7310.n152 3.514
R3269 w_6940_7310.n300 w_6940_7310.n299 3.514
R3270 w_6940_7310.n435 w_6940_7310.n434 3.052
R3271 w_6940_7310.n429 w_6940_7310.n428 3.052
R3272 w_6940_7310.n423 w_6940_7310.n422 3.052
R3273 w_6940_7310.n417 w_6940_7310.n416 3.052
R3274 w_6940_7310.n411 w_6940_7310.n410 3.052
R3275 w_6940_7310.n375 w_6940_7310.n374 3.052
R3276 w_6940_7310.n403 w_6940_7310.n402 3.052
R3277 w_6940_7310.n397 w_6940_7310.n396 3.052
R3278 w_6940_7310.n391 w_6940_7310.n390 3.052
R3279 w_6940_7310.n385 w_6940_7310.n384 3.052
R3280 w_6940_7310.n511 w_6940_7310.n510 3.052
R3281 w_6940_7310.n505 w_6940_7310.n504 3.052
R3282 w_6940_7310.n499 w_6940_7310.n498 3.052
R3283 w_6940_7310.n493 w_6940_7310.n492 3.052
R3284 w_6940_7310.n487 w_6940_7310.n486 3.052
R3285 w_6940_7310.n482 w_6940_7310.n481 3.052
R3286 w_6940_7310.n475 w_6940_7310.n474 3.052
R3287 w_6940_7310.n469 w_6940_7310.n468 3.052
R3288 w_6940_7310.n463 w_6940_7310.n462 3.052
R3289 w_6940_7310.n457 w_6940_7310.n456 3.052
R3290 w_6940_7310.n133 w_6940_7310.n132 3.052
R3291 w_6940_7310.n127 w_6940_7310.n126 3.052
R3292 w_6940_7310.n121 w_6940_7310.n120 3.052
R3293 w_6940_7310.n115 w_6940_7310.n114 3.052
R3294 w_6940_7310.n109 w_6940_7310.n108 3.052
R3295 w_6940_7310.n73 w_6940_7310.n72 3.052
R3296 w_6940_7310.n101 w_6940_7310.n100 3.052
R3297 w_6940_7310.n95 w_6940_7310.n94 3.052
R3298 w_6940_7310.n89 w_6940_7310.n88 3.052
R3299 w_6940_7310.n83 w_6940_7310.n82 3.052
R3300 w_6940_7310.n283 w_6940_7310.n282 3.052
R3301 w_6940_7310.n277 w_6940_7310.n276 3.052
R3302 w_6940_7310.n271 w_6940_7310.n270 3.052
R3303 w_6940_7310.n265 w_6940_7310.n264 3.052
R3304 w_6940_7310.n259 w_6940_7310.n258 3.052
R3305 w_6940_7310.n254 w_6940_7310.n253 3.052
R3306 w_6940_7310.n247 w_6940_7310.n246 3.052
R3307 w_6940_7310.n241 w_6940_7310.n240 3.052
R3308 w_6940_7310.n235 w_6940_7310.n234 3.052
R3309 w_6940_7310.n229 w_6940_7310.n228 3.052
R3310 w_6940_7310.n379 w_6940_7310.n378 2.91
R3311 w_6940_7310.n451 w_6940_7310.n450 2.91
R3312 w_6940_7310.n77 w_6940_7310.n76 2.91
R3313 w_6940_7310.n223 w_6940_7310.n222 2.91
R3314 w_6940_7310.n524 w_6940_7310.n523 2.351
R3315 w_6940_7310.n294 w_6940_7310.n218 0.768
R3316 w_6940_7310.n446 w_6940_7310.n370 0.75
R3317 w_6940_7310.n157 w_6940_7310.n155 0.713
R3318 w_6940_7310.n6 w_6940_7310.n5 0.697
R3319 w_6940_7310.n6 w_6940_7310.n4 0.697
R3320 w_6940_7310.n7 w_6940_7310.n6 0.697
R3321 w_6940_7310.n6 w_6940_7310.n3 0.697
R3322 w_6940_7310.n6 w_6940_7310.n2 0.697
R3323 w_6940_7310.n6 w_6940_7310.n1 0.697
R3324 w_6940_7310.n304 w_6940_7310.n302 0.668
R3325 w_6940_7310.n15 w_6940_7310.n13 0.652
R3326 w_6940_7310.n383 w_6940_7310.n381 0.652
R3327 w_6940_7310.n455 w_6940_7310.n453 0.652
R3328 w_6940_7310.n81 w_6940_7310.n79 0.652
R3329 w_6940_7310.n227 w_6940_7310.n225 0.652
R3330 w_6940_7310.n147 w_6940_7310.n146 0.592
R3331 w_6940_7310.n523 w_6940_7310.n522 0.57
R3332 w_6940_7310.n522 w_6940_7310.n446 0.57
R3333 w_6940_7310.n523 w_6940_7310.n295 0.57
R3334 w_6940_7310.n295 w_6940_7310.n294 0.57
R3335 w_6940_7310.n446 w_6940_7310.n445 0.208
R3336 w_6940_7310.n522 w_6940_7310.n521 0.208
R3337 w_6940_7310.n295 w_6940_7310.n143 0.208
R3338 w_6940_7310.n294 w_6940_7310.n293 0.208
R3339 w_6940_7310.n523 w_6940_7310.n68 0.208
R3340 w_6940_7310.n531 w_6940_7310.n530 0.106
R3341 w_6940_7310.n533 w_6940_7310.n532 0.106
R3342 w_6940_7310.n527 w_6940_7310.n526 0.106
R3343 w_6940_7310.n525 w_6940_7310.n524 0.106
R3344 w_6940_7310.n534 w_6940_7310.n528 0.106
R3345 w_6940_7310.n530 w_6940_7310.n529 0.083
R3346 w_6940_7310.n532 w_6940_7310.n531 0.083
R3347 w_6940_7310.n528 w_6940_7310.n527 0.083
R3348 w_6940_7310.n526 w_6940_7310.n525 0.083
R3349 w_6940_7310.n534 w_6940_7310.n533 0.083
R3350 w_6940_7310.n340 w_6940_7310.n338 0.047
R3351 w_6940_7310.n185 w_6940_7310.n181 0.046
R3352 w_6940_7310.n218 w_6940_7310.n217 0.045
R3353 w_6940_7310.n333 w_6940_7310.n328 0.043
R3354 w_6940_7310.n189 w_6940_7310.n187 0.042
R3355 w_6940_7310.n370 w_6940_7310.n369 0.04
R3356 w_6940_7310.n369 w_6940_7310.n367 0.032
R3357 w_6940_7310.n367 w_6940_7310.n364 0.032
R3358 w_6940_7310.n364 w_6940_7310.n362 0.032
R3359 w_6940_7310.n362 w_6940_7310.n358 0.032
R3360 w_6940_7310.n358 w_6940_7310.n356 0.032
R3361 w_6940_7310.n356 w_6940_7310.n352 0.032
R3362 w_6940_7310.n352 w_6940_7310.n350 0.032
R3363 w_6940_7310.n350 w_6940_7310.n346 0.032
R3364 w_6940_7310.n346 w_6940_7310.n344 0.032
R3365 w_6940_7310.n344 w_6940_7310.n340 0.032
R3366 w_6940_7310.n328 w_6940_7310.n326 0.032
R3367 w_6940_7310.n326 w_6940_7310.n322 0.032
R3368 w_6940_7310.n322 w_6940_7310.n320 0.032
R3369 w_6940_7310.n320 w_6940_7310.n316 0.032
R3370 w_6940_7310.n316 w_6940_7310.n314 0.032
R3371 w_6940_7310.n314 w_6940_7310.n310 0.032
R3372 w_6940_7310.n310 w_6940_7310.n308 0.032
R3373 w_6940_7310.n308 w_6940_7310.n304 0.032
R3374 w_6940_7310.n415 w_6940_7310.n413 0.031
R3375 w_6940_7310.n491 w_6940_7310.n489 0.031
R3376 w_6940_7310.n113 w_6940_7310.n111 0.031
R3377 w_6940_7310.n263 w_6940_7310.n261 0.031
R3378 w_6940_7310.n42 w_6940_7310.n40 0.031
R3379 w_6940_7310.n217 w_6940_7310.n215 0.031
R3380 w_6940_7310.n215 w_6940_7310.n212 0.031
R3381 w_6940_7310.n212 w_6940_7310.n210 0.031
R3382 w_6940_7310.n210 w_6940_7310.n207 0.031
R3383 w_6940_7310.n207 w_6940_7310.n205 0.031
R3384 w_6940_7310.n205 w_6940_7310.n201 0.031
R3385 w_6940_7310.n201 w_6940_7310.n199 0.031
R3386 w_6940_7310.n199 w_6940_7310.n195 0.031
R3387 w_6940_7310.n195 w_6940_7310.n193 0.031
R3388 w_6940_7310.n193 w_6940_7310.n189 0.031
R3389 w_6940_7310.n181 w_6940_7310.n179 0.031
R3390 w_6940_7310.n179 w_6940_7310.n175 0.031
R3391 w_6940_7310.n175 w_6940_7310.n173 0.031
R3392 w_6940_7310.n173 w_6940_7310.n169 0.031
R3393 w_6940_7310.n169 w_6940_7310.n167 0.031
R3394 w_6940_7310.n167 w_6940_7310.n163 0.031
R3395 w_6940_7310.n163 w_6940_7310.n161 0.031
R3396 w_6940_7310.n161 w_6940_7310.n157 0.031
R3397 w_6940_7310.n338 w_6940_7310.n334 0.031
R3398 w_6940_7310.n186 w_6940_7310.n185 0.03
R3399 w_6940_7310.n408 w_6940_7310.n407 0.029
R3400 w_6940_7310.n484 w_6940_7310.n479 0.029
R3401 w_6940_7310.n106 w_6940_7310.n105 0.029
R3402 w_6940_7310.n256 w_6940_7310.n251 0.029
R3403 w_6940_7310.n36 w_6940_7310.n35 0.029
R3404 w_6940_7310.n445 w_6940_7310.n444 0.027
R3405 w_6940_7310.n521 w_6940_7310.n520 0.027
R3406 w_6940_7310.n143 w_6940_7310.n142 0.027
R3407 w_6940_7310.n293 w_6940_7310.n292 0.027
R3408 w_6940_7310.n68 w_6940_7310.n67 0.027
R3409 w_6940_7310.n444 w_6940_7310.n442 0.021
R3410 w_6940_7310.n442 w_6940_7310.n439 0.021
R3411 w_6940_7310.n439 w_6940_7310.n437 0.021
R3412 w_6940_7310.n437 w_6940_7310.n433 0.021
R3413 w_6940_7310.n433 w_6940_7310.n431 0.021
R3414 w_6940_7310.n431 w_6940_7310.n427 0.021
R3415 w_6940_7310.n427 w_6940_7310.n425 0.021
R3416 w_6940_7310.n425 w_6940_7310.n421 0.021
R3417 w_6940_7310.n421 w_6940_7310.n419 0.021
R3418 w_6940_7310.n419 w_6940_7310.n415 0.021
R3419 w_6940_7310.n407 w_6940_7310.n405 0.021
R3420 w_6940_7310.n405 w_6940_7310.n401 0.021
R3421 w_6940_7310.n401 w_6940_7310.n399 0.021
R3422 w_6940_7310.n399 w_6940_7310.n395 0.021
R3423 w_6940_7310.n395 w_6940_7310.n393 0.021
R3424 w_6940_7310.n393 w_6940_7310.n389 0.021
R3425 w_6940_7310.n389 w_6940_7310.n387 0.021
R3426 w_6940_7310.n387 w_6940_7310.n383 0.021
R3427 w_6940_7310.n520 w_6940_7310.n518 0.021
R3428 w_6940_7310.n518 w_6940_7310.n515 0.021
R3429 w_6940_7310.n515 w_6940_7310.n513 0.021
R3430 w_6940_7310.n513 w_6940_7310.n509 0.021
R3431 w_6940_7310.n509 w_6940_7310.n507 0.021
R3432 w_6940_7310.n507 w_6940_7310.n503 0.021
R3433 w_6940_7310.n503 w_6940_7310.n501 0.021
R3434 w_6940_7310.n501 w_6940_7310.n497 0.021
R3435 w_6940_7310.n497 w_6940_7310.n495 0.021
R3436 w_6940_7310.n495 w_6940_7310.n491 0.021
R3437 w_6940_7310.n479 w_6940_7310.n477 0.021
R3438 w_6940_7310.n477 w_6940_7310.n473 0.021
R3439 w_6940_7310.n473 w_6940_7310.n471 0.021
R3440 w_6940_7310.n471 w_6940_7310.n467 0.021
R3441 w_6940_7310.n467 w_6940_7310.n465 0.021
R3442 w_6940_7310.n465 w_6940_7310.n461 0.021
R3443 w_6940_7310.n461 w_6940_7310.n459 0.021
R3444 w_6940_7310.n459 w_6940_7310.n455 0.021
R3445 w_6940_7310.n142 w_6940_7310.n140 0.021
R3446 w_6940_7310.n140 w_6940_7310.n137 0.021
R3447 w_6940_7310.n137 w_6940_7310.n135 0.021
R3448 w_6940_7310.n135 w_6940_7310.n131 0.021
R3449 w_6940_7310.n131 w_6940_7310.n129 0.021
R3450 w_6940_7310.n129 w_6940_7310.n125 0.021
R3451 w_6940_7310.n125 w_6940_7310.n123 0.021
R3452 w_6940_7310.n123 w_6940_7310.n119 0.021
R3453 w_6940_7310.n119 w_6940_7310.n117 0.021
R3454 w_6940_7310.n117 w_6940_7310.n113 0.021
R3455 w_6940_7310.n105 w_6940_7310.n103 0.021
R3456 w_6940_7310.n103 w_6940_7310.n99 0.021
R3457 w_6940_7310.n99 w_6940_7310.n97 0.021
R3458 w_6940_7310.n97 w_6940_7310.n93 0.021
R3459 w_6940_7310.n93 w_6940_7310.n91 0.021
R3460 w_6940_7310.n91 w_6940_7310.n87 0.021
R3461 w_6940_7310.n87 w_6940_7310.n85 0.021
R3462 w_6940_7310.n85 w_6940_7310.n81 0.021
R3463 w_6940_7310.n292 w_6940_7310.n290 0.021
R3464 w_6940_7310.n290 w_6940_7310.n287 0.021
R3465 w_6940_7310.n287 w_6940_7310.n285 0.021
R3466 w_6940_7310.n285 w_6940_7310.n281 0.021
R3467 w_6940_7310.n281 w_6940_7310.n279 0.021
R3468 w_6940_7310.n279 w_6940_7310.n275 0.021
R3469 w_6940_7310.n275 w_6940_7310.n273 0.021
R3470 w_6940_7310.n273 w_6940_7310.n269 0.021
R3471 w_6940_7310.n269 w_6940_7310.n267 0.021
R3472 w_6940_7310.n267 w_6940_7310.n263 0.021
R3473 w_6940_7310.n251 w_6940_7310.n249 0.021
R3474 w_6940_7310.n249 w_6940_7310.n245 0.021
R3475 w_6940_7310.n245 w_6940_7310.n243 0.021
R3476 w_6940_7310.n243 w_6940_7310.n239 0.021
R3477 w_6940_7310.n239 w_6940_7310.n237 0.021
R3478 w_6940_7310.n237 w_6940_7310.n233 0.021
R3479 w_6940_7310.n233 w_6940_7310.n231 0.021
R3480 w_6940_7310.n231 w_6940_7310.n227 0.021
R3481 w_6940_7310.n67 w_6940_7310.n65 0.021
R3482 w_6940_7310.n65 w_6940_7310.n62 0.021
R3483 w_6940_7310.n62 w_6940_7310.n60 0.021
R3484 w_6940_7310.n60 w_6940_7310.n57 0.021
R3485 w_6940_7310.n57 w_6940_7310.n55 0.021
R3486 w_6940_7310.n55 w_6940_7310.n52 0.021
R3487 w_6940_7310.n52 w_6940_7310.n50 0.021
R3488 w_6940_7310.n50 w_6940_7310.n47 0.021
R3489 w_6940_7310.n47 w_6940_7310.n45 0.021
R3490 w_6940_7310.n45 w_6940_7310.n42 0.021
R3491 w_6940_7310.n35 w_6940_7310.n33 0.021
R3492 w_6940_7310.n33 w_6940_7310.n30 0.021
R3493 w_6940_7310.n30 w_6940_7310.n28 0.021
R3494 w_6940_7310.n28 w_6940_7310.n25 0.021
R3495 w_6940_7310.n25 w_6940_7310.n23 0.021
R3496 w_6940_7310.n23 w_6940_7310.n20 0.021
R3497 w_6940_7310.n20 w_6940_7310.n18 0.021
R3498 w_6940_7310.n18 w_6940_7310.n15 0.021
R3499 w_6940_7310.n413 w_6940_7310.n409 0.021
R3500 w_6940_7310.n489 w_6940_7310.n485 0.021
R3501 w_6940_7310.n111 w_6940_7310.n107 0.021
R3502 w_6940_7310.n261 w_6940_7310.n257 0.021
R3503 w_6940_7310.n40 w_6940_7310.n37 0.021
R3504 w_6940_7310.n334 w_6940_7310.n333 0.009
R3505 w_6940_7310.n187 w_6940_7310.n186 0.009
R3506 w_6940_7310.n409 w_6940_7310.n408 0.006
R3507 w_6940_7310.n485 w_6940_7310.n484 0.006
R3508 w_6940_7310.n107 w_6940_7310.n106 0.006
R3509 w_6940_7310.n257 w_6940_7310.n256 0.006
R3510 w_6940_7310.n37 w_6940_7310.n36 0.006
R3511 a_7170_7410.n7 a_7170_7410.t14 708.072
R3512 a_7170_7410.n9 a_7170_7410.t16 708.056
R3513 a_7170_7410.n11 a_7170_7410.t17 708.054
R3514 a_7170_7410.n11 a_7170_7410.t15 708.054
R3515 a_7170_7410.n9 a_7170_7410.t20 708.05
R3516 a_7170_7410.n7 a_7170_7410.t22 708.038
R3517 a_7170_7410.n6 a_7170_7410.t23 388.574
R3518 a_7170_7410.n6 a_7170_7410.t21 388.524
R3519 a_7170_7410.n12 a_7170_7410.t19 388.509
R3520 a_7170_7410.n12 a_7170_7410.t24 388.509
R3521 a_7170_7410.n10 a_7170_7410.t13 388.509
R3522 a_7170_7410.n10 a_7170_7410.t18 388.509
R3523 a_7170_7410.n13 a_7170_7410.t1 5.713
R3524 a_7170_7410.n13 a_7170_7410.t7 5.713
R3525 a_7170_7410.n5 a_7170_7410.t2 5.713
R3526 a_7170_7410.n5 a_7170_7410.t8 5.713
R3527 a_7170_7410.n3 a_7170_7410.t4 5.713
R3528 a_7170_7410.n3 a_7170_7410.t11 5.713
R3529 a_7170_7410.n4 a_7170_7410.t6 3.48
R3530 a_7170_7410.n4 a_7170_7410.t3 3.48
R3531 a_7170_7410.n2 a_7170_7410.t9 3.48
R3532 a_7170_7410.n2 a_7170_7410.t10 3.48
R3533 a_7170_7410.n14 a_7170_7410.t5 3.48
R3534 a_7170_7410.t0 a_7170_7410.n14 3.48
R3535 a_7170_7410.t12 a_7170_7410.n1 2.751
R3536 a_7170_7410.n1 a_7170_7410.n11 2.272
R3537 a_7170_7410.n8 a_7170_7410.n7 2.265
R3538 a_7170_7410.n0 a_7170_7410.n9 2.178
R3539 a_7170_7410.n5 a_7170_7410.n4 1.164
R3540 a_7170_7410.n3 a_7170_7410.n2 1.164
R3541 a_7170_7410.n14 a_7170_7410.n13 1.112
R3542 a_7170_7410.n1 a_7170_7410.n0 0.841
R3543 a_7170_7410.n0 a_7170_7410.n8 0.804
R3544 a_7170_7410.n8 a_7170_7410.n6 0.328
R3545 a_7170_7410.n1 a_7170_7410.n12 0.29
R3546 a_7170_7410.t12 a_7170_7410.n3 0.2
R3547 a_7170_7410.t12 a_7170_7410.n5 0.2
R3548 a_7170_7410.n13 a_7170_7410.t12 0.2
R3549 a_7170_7410.n0 a_7170_7410.n10 0.162
R3550 a_7100_7313.n7 a_7100_7313.t14 708.034
R3551 a_7100_7313.n6 a_7100_7313.t15 708.034
R3552 a_7100_7313.n9 a_7100_7313.t16 708.034
R3553 a_7100_7313.n7 a_7100_7313.t24 708.034
R3554 a_7100_7313.n6 a_7100_7313.t21 708.034
R3555 a_7100_7313.n9 a_7100_7313.t23 708.034
R3556 a_7100_7313.n10 a_7100_7313.t18 388.664
R3557 a_7100_7313.n8 a_7100_7313.t13 388.587
R3558 a_7100_7313.n8 a_7100_7313.t20 388.587
R3559 a_7100_7313.n5 a_7100_7313.t17 388.587
R3560 a_7100_7313.n5 a_7100_7313.t12 388.587
R3561 a_7100_7313.n10 a_7100_7313.t22 388.543
R3562 a_7100_7313.n18 a_7100_7313.t1 5.713
R3563 a_7100_7313.n18 a_7100_7313.t2 5.713
R3564 a_7100_7313.n14 a_7100_7313.t4 5.713
R3565 a_7100_7313.n14 a_7100_7313.t5 5.713
R3566 a_7100_7313.n3 a_7100_7313.t0 5.713
R3567 a_7100_7313.n3 a_7100_7313.t3 5.713
R3568 a_7100_7313.n13 a_7100_7313.t7 3.48
R3569 a_7100_7313.n13 a_7100_7313.t9 3.48
R3570 a_7100_7313.n2 a_7100_7313.t8 3.48
R3571 a_7100_7313.n2 a_7100_7313.t10 3.48
R3572 a_7100_7313.n20 a_7100_7313.t6 3.48
R3573 a_7100_7313.t11 a_7100_7313.n20 3.48
R3574 a_7100_7313.n12 a_7100_7313.n0 2.556
R3575 a_7100_7313.n0 a_7100_7313.n6 2.489
R3576 a_7100_7313.n11 a_7100_7313.n9 2.478
R3577 a_7100_7313.n1 a_7100_7313.n7 2.348
R3578 a_7100_7313.n0 a_7100_7313.n1 0.841
R3579 a_7100_7313.n1 a_7100_7313.n11 0.819
R3580 a_7100_7313.n15 a_7100_7313.n13 0.701
R3581 a_7100_7313.n4 a_7100_7313.n2 0.701
R3582 a_7100_7313.n20 a_7100_7313.n19 0.701
R3583 a_7100_7313.n15 a_7100_7313.n14 0.463
R3584 a_7100_7313.n4 a_7100_7313.n3 0.463
R3585 a_7100_7313.n19 a_7100_7313.n18 0.419
R3586 a_7100_7313.t19 a_7100_7313.n4 0.141
R3587 a_7100_7313.n17 a_7100_7313.n16 0.135
R3588 a_7100_7313.n16 a_7100_7313.n15 0.116
R3589 a_7100_7313.n19 a_7100_7313.n17 0.112
R3590 a_7100_7313.n11 a_7100_7313.n10 0.099
R3591 a_7100_7313.n0 a_7100_7313.n5 0.077
R3592 a_7100_7313.n17 a_7100_7313.n12 0.058
R3593 a_7100_7313.n1 a_7100_7313.n8 0.03
R3594 a_7100_7313.n12 a_7100_7313.t19 0.025
R3595 w_19680_7310.n293 w_19680_7310.t10 112.822
R3596 w_19680_7310.n368 w_19680_7310.t14 112.822
R3597 w_19680_7310.n368 w_19680_7310.t22 112.822
R3598 w_19680_7310.n444 w_19680_7310.t28 112.822
R3599 w_19680_7310.n444 w_19680_7310.t12 112.822
R3600 w_19680_7310.n0 w_19680_7310.t16 112.822
R3601 w_19680_7310.n0 w_19680_7310.t18 112.822
R3602 w_19680_7310.n196 w_19680_7310.t20 112.822
R3603 w_19680_7310.n196 w_19680_7310.t6 112.822
R3604 w_19680_7310.n147 w_19680_7310.t8 112.822
R3605 w_19680_7310.n147 w_19680_7310.t24 112.822
R3606 w_19680_7310.n42 w_19680_7310.t26 112.822
R3607 w_19680_7310.n203 w_19680_7310.n200 20.092
R3608 w_19680_7310.n261 w_19680_7310.n260 16.607
R3609 w_19680_7310.n115 w_19680_7310.n114 16.289
R3610 w_19680_7310.n412 w_19680_7310.n411 16.289
R3611 w_19680_7310.n336 w_19680_7310.n335 16.289
R3612 w_19680_7310.n500 w_19680_7310.n499 16.288
R3613 w_19680_7310.n50 w_19680_7310.n46 12.923
R3614 w_19680_7310.n266 w_19680_7310.n262 12.641
R3615 w_19680_7310.n8 w_19680_7310.n4 12.629
R3616 w_19680_7310.n341 w_19680_7310.n337 12.629
R3617 w_19680_7310.n417 w_19680_7310.n413 12.629
R3618 w_19680_7310.n120 w_19680_7310.n116 12.629
R3619 w_19680_7310.n40 w_19680_7310.n39 12.369
R3620 w_19680_7310.n268 w_19680_7310.n267 9.3
R3621 w_19680_7310.n274 w_19680_7310.n273 9.3
R3622 w_19680_7310.n280 w_19680_7310.n279 9.3
R3623 w_19680_7310.n286 w_19680_7310.n285 9.3
R3624 w_19680_7310.n292 w_19680_7310.n291 9.3
R3625 w_19680_7310.n304 w_19680_7310.n303 9.3
R3626 w_19680_7310.n310 w_19680_7310.n309 9.3
R3627 w_19680_7310.n316 w_19680_7310.n315 9.3
R3628 w_19680_7310.n322 w_19680_7310.n321 9.3
R3629 w_19680_7310.n328 w_19680_7310.n327 9.3
R3630 w_19680_7310.n333 w_19680_7310.n332 9.3
R3631 w_19680_7310.n343 w_19680_7310.n342 9.3
R3632 w_19680_7310.n349 w_19680_7310.n348 9.3
R3633 w_19680_7310.n355 w_19680_7310.n354 9.3
R3634 w_19680_7310.n361 w_19680_7310.n360 9.3
R3635 w_19680_7310.n367 w_19680_7310.n366 9.3
R3636 w_19680_7310.n379 w_19680_7310.n378 9.3
R3637 w_19680_7310.n385 w_19680_7310.n384 9.3
R3638 w_19680_7310.n391 w_19680_7310.n390 9.3
R3639 w_19680_7310.n397 w_19680_7310.n396 9.3
R3640 w_19680_7310.n403 w_19680_7310.n402 9.3
R3641 w_19680_7310.n408 w_19680_7310.n407 9.3
R3642 w_19680_7310.n419 w_19680_7310.n418 9.3
R3643 w_19680_7310.n425 w_19680_7310.n424 9.3
R3644 w_19680_7310.n431 w_19680_7310.n430 9.3
R3645 w_19680_7310.n437 w_19680_7310.n436 9.3
R3646 w_19680_7310.n443 w_19680_7310.n442 9.3
R3647 w_19680_7310.n455 w_19680_7310.n454 9.3
R3648 w_19680_7310.n461 w_19680_7310.n460 9.3
R3649 w_19680_7310.n467 w_19680_7310.n466 9.3
R3650 w_19680_7310.n473 w_19680_7310.n472 9.3
R3651 w_19680_7310.n479 w_19680_7310.n478 9.3
R3652 w_19680_7310.n484 w_19680_7310.n483 9.3
R3653 w_19680_7310.n112 w_19680_7310.n111 9.3
R3654 w_19680_7310.n52 w_19680_7310.n51 9.3
R3655 w_19680_7310.n58 w_19680_7310.n57 9.3
R3656 w_19680_7310.n64 w_19680_7310.n63 9.3
R3657 w_19680_7310.n70 w_19680_7310.n69 9.3
R3658 w_19680_7310.n76 w_19680_7310.n75 9.3
R3659 w_19680_7310.n84 w_19680_7310.n83 9.3
R3660 w_19680_7310.n90 w_19680_7310.n89 9.3
R3661 w_19680_7310.n96 w_19680_7310.n95 9.3
R3662 w_19680_7310.n102 w_19680_7310.n101 9.3
R3663 w_19680_7310.n107 w_19680_7310.n106 9.3
R3664 w_19680_7310.n122 w_19680_7310.n121 9.3
R3665 w_19680_7310.n128 w_19680_7310.n127 9.3
R3666 w_19680_7310.n134 w_19680_7310.n133 9.3
R3667 w_19680_7310.n140 w_19680_7310.n139 9.3
R3668 w_19680_7310.n146 w_19680_7310.n145 9.3
R3669 w_19680_7310.n158 w_19680_7310.n157 9.3
R3670 w_19680_7310.n164 w_19680_7310.n163 9.3
R3671 w_19680_7310.n170 w_19680_7310.n169 9.3
R3672 w_19680_7310.n176 w_19680_7310.n175 9.3
R3673 w_19680_7310.n182 w_19680_7310.n181 9.3
R3674 w_19680_7310.n187 w_19680_7310.n186 9.3
R3675 w_19680_7310.n126 w_19680_7310.n125 9.3
R3676 w_19680_7310.n132 w_19680_7310.n131 9.3
R3677 w_19680_7310.n138 w_19680_7310.n137 9.3
R3678 w_19680_7310.n144 w_19680_7310.n143 9.3
R3679 w_19680_7310.n162 w_19680_7310.n161 9.3
R3680 w_19680_7310.n168 w_19680_7310.n167 9.3
R3681 w_19680_7310.n174 w_19680_7310.n173 9.3
R3682 w_19680_7310.n180 w_19680_7310.n179 9.3
R3683 w_19680_7310.n185 w_19680_7310.n184 9.3
R3684 w_19680_7310.n423 w_19680_7310.n422 9.3
R3685 w_19680_7310.n429 w_19680_7310.n428 9.3
R3686 w_19680_7310.n435 w_19680_7310.n434 9.3
R3687 w_19680_7310.n441 w_19680_7310.n440 9.3
R3688 w_19680_7310.n459 w_19680_7310.n458 9.3
R3689 w_19680_7310.n465 w_19680_7310.n464 9.3
R3690 w_19680_7310.n471 w_19680_7310.n470 9.3
R3691 w_19680_7310.n477 w_19680_7310.n476 9.3
R3692 w_19680_7310.n482 w_19680_7310.n481 9.3
R3693 w_19680_7310.n347 w_19680_7310.n346 9.3
R3694 w_19680_7310.n353 w_19680_7310.n352 9.3
R3695 w_19680_7310.n359 w_19680_7310.n358 9.3
R3696 w_19680_7310.n365 w_19680_7310.n364 9.3
R3697 w_19680_7310.n383 w_19680_7310.n382 9.3
R3698 w_19680_7310.n389 w_19680_7310.n388 9.3
R3699 w_19680_7310.n395 w_19680_7310.n394 9.3
R3700 w_19680_7310.n401 w_19680_7310.n400 9.3
R3701 w_19680_7310.n406 w_19680_7310.n405 9.3
R3702 w_19680_7310.n272 w_19680_7310.n271 9.3
R3703 w_19680_7310.n278 w_19680_7310.n277 9.3
R3704 w_19680_7310.n284 w_19680_7310.n283 9.3
R3705 w_19680_7310.n290 w_19680_7310.n289 9.3
R3706 w_19680_7310.n308 w_19680_7310.n307 9.3
R3707 w_19680_7310.n314 w_19680_7310.n313 9.3
R3708 w_19680_7310.n320 w_19680_7310.n319 9.3
R3709 w_19680_7310.n326 w_19680_7310.n325 9.3
R3710 w_19680_7310.n331 w_19680_7310.n330 9.3
R3711 w_19680_7310.n56 w_19680_7310.n55 9.3
R3712 w_19680_7310.n62 w_19680_7310.n61 9.3
R3713 w_19680_7310.n68 w_19680_7310.n67 9.3
R3714 w_19680_7310.n74 w_19680_7310.n73 9.3
R3715 w_19680_7310.n88 w_19680_7310.n87 9.3
R3716 w_19680_7310.n94 w_19680_7310.n93 9.3
R3717 w_19680_7310.n100 w_19680_7310.n99 9.3
R3718 w_19680_7310.n105 w_19680_7310.n104 9.3
R3719 w_19680_7310.n110 w_19680_7310.n109 9.3
R3720 w_19680_7310.n205 w_19680_7310.n204 9.3
R3721 w_19680_7310.n208 w_19680_7310.n207 9.3
R3722 w_19680_7310.n210 w_19680_7310.n209 9.3
R3723 w_19680_7310.n213 w_19680_7310.n212 9.3
R3724 w_19680_7310.n215 w_19680_7310.n214 9.3
R3725 w_19680_7310.n218 w_19680_7310.n217 9.3
R3726 w_19680_7310.n220 w_19680_7310.n219 9.3
R3727 w_19680_7310.n223 w_19680_7310.n222 9.3
R3728 w_19680_7310.n225 w_19680_7310.n224 9.3
R3729 w_19680_7310.n232 w_19680_7310.n231 9.3
R3730 w_19680_7310.n235 w_19680_7310.n234 9.3
R3731 w_19680_7310.n237 w_19680_7310.n236 9.3
R3732 w_19680_7310.n240 w_19680_7310.n239 9.3
R3733 w_19680_7310.n242 w_19680_7310.n241 9.3
R3734 w_19680_7310.n245 w_19680_7310.n244 9.3
R3735 w_19680_7310.n247 w_19680_7310.n246 9.3
R3736 w_19680_7310.n250 w_19680_7310.n249 9.3
R3737 w_19680_7310.n252 w_19680_7310.n251 9.3
R3738 w_19680_7310.n255 w_19680_7310.n254 9.3
R3739 w_19680_7310.n257 w_19680_7310.n256 9.3
R3740 w_19680_7310.n10 w_19680_7310.n9 9.3
R3741 w_19680_7310.n14 w_19680_7310.n13 9.3
R3742 w_19680_7310.n16 w_19680_7310.n15 9.3
R3743 w_19680_7310.n20 w_19680_7310.n19 9.3
R3744 w_19680_7310.n22 w_19680_7310.n21 9.3
R3745 w_19680_7310.n26 w_19680_7310.n25 9.3
R3746 w_19680_7310.n28 w_19680_7310.n27 9.3
R3747 w_19680_7310.n32 w_19680_7310.n31 9.3
R3748 w_19680_7310.n34 w_19680_7310.n33 9.3
R3749 w_19680_7310.n532 w_19680_7310.n531 9.3
R3750 w_19680_7310.n530 w_19680_7310.n529 9.3
R3751 w_19680_7310.n526 w_19680_7310.n525 9.3
R3752 w_19680_7310.n524 w_19680_7310.n523 9.3
R3753 w_19680_7310.n520 w_19680_7310.n519 9.3
R3754 w_19680_7310.n518 w_19680_7310.n517 9.3
R3755 w_19680_7310.n514 w_19680_7310.n513 9.3
R3756 w_19680_7310.n512 w_19680_7310.n511 9.3
R3757 w_19680_7310.n508 w_19680_7310.n507 9.3
R3758 w_19680_7310.n506 w_19680_7310.n505 9.3
R3759 w_19680_7310.n503 w_19680_7310.n502 9.3
R3760 w_19680_7310.n119 w_19680_7310.n118 8.855
R3761 w_19680_7310.n125 w_19680_7310.n124 8.855
R3762 w_19680_7310.n131 w_19680_7310.n130 8.855
R3763 w_19680_7310.n137 w_19680_7310.n136 8.855
R3764 w_19680_7310.n143 w_19680_7310.n142 8.855
R3765 w_19680_7310.n150 w_19680_7310.n149 8.855
R3766 w_19680_7310.n155 w_19680_7310.n154 8.855
R3767 w_19680_7310.n161 w_19680_7310.n160 8.855
R3768 w_19680_7310.n167 w_19680_7310.n166 8.855
R3769 w_19680_7310.n173 w_19680_7310.n172 8.855
R3770 w_19680_7310.n179 w_19680_7310.n178 8.855
R3771 w_19680_7310.n184 w_19680_7310.n183 8.855
R3772 w_19680_7310.n7 w_19680_7310.n6 8.855
R3773 w_19680_7310.n416 w_19680_7310.n415 8.855
R3774 w_19680_7310.n422 w_19680_7310.n421 8.855
R3775 w_19680_7310.n428 w_19680_7310.n427 8.855
R3776 w_19680_7310.n434 w_19680_7310.n433 8.855
R3777 w_19680_7310.n440 w_19680_7310.n439 8.855
R3778 w_19680_7310.n447 w_19680_7310.n446 8.855
R3779 w_19680_7310.n452 w_19680_7310.n451 8.855
R3780 w_19680_7310.n458 w_19680_7310.n457 8.855
R3781 w_19680_7310.n464 w_19680_7310.n463 8.855
R3782 w_19680_7310.n470 w_19680_7310.n469 8.855
R3783 w_19680_7310.n476 w_19680_7310.n475 8.855
R3784 w_19680_7310.n481 w_19680_7310.n480 8.855
R3785 w_19680_7310.n340 w_19680_7310.n339 8.855
R3786 w_19680_7310.n346 w_19680_7310.n345 8.855
R3787 w_19680_7310.n352 w_19680_7310.n351 8.855
R3788 w_19680_7310.n358 w_19680_7310.n357 8.855
R3789 w_19680_7310.n364 w_19680_7310.n363 8.855
R3790 w_19680_7310.n371 w_19680_7310.n370 8.855
R3791 w_19680_7310.n376 w_19680_7310.n375 8.855
R3792 w_19680_7310.n382 w_19680_7310.n381 8.855
R3793 w_19680_7310.n388 w_19680_7310.n387 8.855
R3794 w_19680_7310.n394 w_19680_7310.n393 8.855
R3795 w_19680_7310.n400 w_19680_7310.n399 8.855
R3796 w_19680_7310.n405 w_19680_7310.n404 8.855
R3797 w_19680_7310.n265 w_19680_7310.n264 8.855
R3798 w_19680_7310.n271 w_19680_7310.n270 8.855
R3799 w_19680_7310.n277 w_19680_7310.n276 8.855
R3800 w_19680_7310.n283 w_19680_7310.n282 8.855
R3801 w_19680_7310.n289 w_19680_7310.n288 8.855
R3802 w_19680_7310.n296 w_19680_7310.n295 8.855
R3803 w_19680_7310.n301 w_19680_7310.n300 8.855
R3804 w_19680_7310.n307 w_19680_7310.n306 8.855
R3805 w_19680_7310.n313 w_19680_7310.n312 8.855
R3806 w_19680_7310.n319 w_19680_7310.n318 8.855
R3807 w_19680_7310.n325 w_19680_7310.n324 8.855
R3808 w_19680_7310.n330 w_19680_7310.n329 8.855
R3809 w_19680_7310.n49 w_19680_7310.n48 8.855
R3810 w_19680_7310.n55 w_19680_7310.n54 8.855
R3811 w_19680_7310.n61 w_19680_7310.n60 8.855
R3812 w_19680_7310.n67 w_19680_7310.n66 8.855
R3813 w_19680_7310.n73 w_19680_7310.n72 8.855
R3814 w_19680_7310.n79 w_19680_7310.n78 8.855
R3815 w_19680_7310.n45 w_19680_7310.n44 8.855
R3816 w_19680_7310.n87 w_19680_7310.n86 8.855
R3817 w_19680_7310.n93 w_19680_7310.n92 8.855
R3818 w_19680_7310.n99 w_19680_7310.n98 8.855
R3819 w_19680_7310.n104 w_19680_7310.n103 8.855
R3820 w_19680_7310.n109 w_19680_7310.n108 8.855
R3821 w_19680_7310.n202 w_19680_7310.n201 8.855
R3822 w_19680_7310.n207 w_19680_7310.n206 8.855
R3823 w_19680_7310.n212 w_19680_7310.n211 8.855
R3824 w_19680_7310.n217 w_19680_7310.n216 8.855
R3825 w_19680_7310.n222 w_19680_7310.n221 8.855
R3826 w_19680_7310.n199 w_19680_7310.n198 8.855
R3827 w_19680_7310.n229 w_19680_7310.n228 8.855
R3828 w_19680_7310.n234 w_19680_7310.n233 8.855
R3829 w_19680_7310.n239 w_19680_7310.n238 8.855
R3830 w_19680_7310.n244 w_19680_7310.n243 8.855
R3831 w_19680_7310.n249 w_19680_7310.n248 8.855
R3832 w_19680_7310.n254 w_19680_7310.n253 8.855
R3833 w_19680_7310.n13 w_19680_7310.n12 8.855
R3834 w_19680_7310.n19 w_19680_7310.n18 8.855
R3835 w_19680_7310.n25 w_19680_7310.n24 8.855
R3836 w_19680_7310.n31 w_19680_7310.n30 8.855
R3837 w_19680_7310.n3 w_19680_7310.n2 8.855
R3838 w_19680_7310.n38 w_19680_7310.n37 8.855
R3839 w_19680_7310.n529 w_19680_7310.n528 8.855
R3840 w_19680_7310.n523 w_19680_7310.n522 8.855
R3841 w_19680_7310.n517 w_19680_7310.n516 8.855
R3842 w_19680_7310.n511 w_19680_7310.n510 8.855
R3843 w_19680_7310.n505 w_19680_7310.n504 8.855
R3844 w_19680_7310.n198 w_19680_7310.n197 7.463
R3845 w_19680_7310.n188 w_19680_7310.n115 6.209
R3846 w_19680_7310.n485 w_19680_7310.n412 6.209
R3847 w_19680_7310.n409 w_19680_7310.n336 6.209
R3848 w_19680_7310.n258 w_19680_7310.n190 6.209
R3849 w_19680_7310.n501 w_19680_7310.n500 6.209
R3850 w_19680_7310.n334 w_19680_7310.n261 6.208
R3851 w_19680_7310.n148 w_19680_7310.n147 5.95
R3852 w_19680_7310.n445 w_19680_7310.n444 5.95
R3853 w_19680_7310.n369 w_19680_7310.n368 5.95
R3854 w_19680_7310.n1 w_19680_7310.n0 5.95
R3855 w_19680_7310.n156 w_19680_7310.n155 5.876
R3856 w_19680_7310.n453 w_19680_7310.n452 5.876
R3857 w_19680_7310.n377 w_19680_7310.n376 5.876
R3858 w_19680_7310.n230 w_19680_7310.n229 5.876
R3859 w_19680_7310.n533 w_19680_7310.n38 5.876
R3860 w_19680_7310.n80 w_19680_7310.n79 5.873
R3861 w_19680_7310.n302 w_19680_7310.n301 5.873
R3862 w_19680_7310.n534 w_19680_7310.t19 5.713
R3863 w_19680_7310.n227 w_19680_7310.t21 5.713
R3864 w_19680_7310.n373 w_19680_7310.t15 5.713
R3865 w_19680_7310.n373 w_19680_7310.t23 5.713
R3866 w_19680_7310.n298 w_19680_7310.t11 5.713
R3867 w_19680_7310.n449 w_19680_7310.t29 5.713
R3868 w_19680_7310.n449 w_19680_7310.t13 5.713
R3869 w_19680_7310.n152 w_19680_7310.t9 5.713
R3870 w_19680_7310.n152 w_19680_7310.t25 5.713
R3871 w_19680_7310.n81 w_19680_7310.t27 5.713
R3872 w_19680_7310.n227 w_19680_7310.t7 5.713
R3873 w_19680_7310.t17 w_19680_7310.n534 5.713
R3874 w_19680_7310.n113 w_19680_7310.n40 5.637
R3875 w_19680_7310.n120 w_19680_7310.n119 5.614
R3876 w_19680_7310.n417 w_19680_7310.n416 5.614
R3877 w_19680_7310.n341 w_19680_7310.n340 5.614
R3878 w_19680_7310.n203 w_19680_7310.n202 5.614
R3879 w_19680_7310.n8 w_19680_7310.n7 5.614
R3880 w_19680_7310.n266 w_19680_7310.n265 5.611
R3881 w_19680_7310.n50 w_19680_7310.n49 5.571
R3882 w_19680_7310.n294 w_19680_7310.n293 5.347
R3883 w_19680_7310.n43 w_19680_7310.n42 5.347
R3884 w_19680_7310.n487 w_19680_7310.t30 4.439
R3885 w_19680_7310.n487 w_19680_7310.t34 4.386
R3886 w_19680_7310.n488 w_19680_7310.t2 4.386
R3887 w_19680_7310.n489 w_19680_7310.t5 4.386
R3888 w_19680_7310.n490 w_19680_7310.t32 4.386
R3889 w_19680_7310.n491 w_19680_7310.t33 4.386
R3890 w_19680_7310.n492 w_19680_7310.t1 4.386
R3891 w_19680_7310.n493 w_19680_7310.t4 4.386
R3892 w_19680_7310.n494 w_19680_7310.t31 4.386
R3893 w_19680_7310.n495 w_19680_7310.t35 4.386
R3894 w_19680_7310.n496 w_19680_7310.t0 4.386
R3895 w_19680_7310.n497 w_19680_7310.t3 4.386
R3896 w_19680_7310.n372 w_19680_7310.n371 4.27
R3897 w_19680_7310.n448 w_19680_7310.n447 4.27
R3898 w_19680_7310.n151 w_19680_7310.n150 4.27
R3899 w_19680_7310.n226 w_19680_7310.n199 4.27
R3900 w_19680_7310.n35 w_19680_7310.n3 4.27
R3901 w_19680_7310.n297 w_19680_7310.n296 4.269
R3902 w_19680_7310.n82 w_19680_7310.n45 4.269
R3903 w_19680_7310.n498 w_19680_7310.n497 3.948
R3904 w_19680_7310.n98 w_19680_7310.n97 3.685
R3905 w_19680_7310.n92 w_19680_7310.n91 3.685
R3906 w_19680_7310.n86 w_19680_7310.n85 3.685
R3907 w_19680_7310.n44 w_19680_7310.n43 3.685
R3908 w_19680_7310.n78 w_19680_7310.n77 3.685
R3909 w_19680_7310.n72 w_19680_7310.n71 3.685
R3910 w_19680_7310.n66 w_19680_7310.n65 3.685
R3911 w_19680_7310.n60 w_19680_7310.n59 3.685
R3912 w_19680_7310.n54 w_19680_7310.n53 3.685
R3913 w_19680_7310.n324 w_19680_7310.n323 3.685
R3914 w_19680_7310.n318 w_19680_7310.n317 3.685
R3915 w_19680_7310.n312 w_19680_7310.n311 3.685
R3916 w_19680_7310.n306 w_19680_7310.n305 3.685
R3917 w_19680_7310.n300 w_19680_7310.n299 3.685
R3918 w_19680_7310.n295 w_19680_7310.n294 3.685
R3919 w_19680_7310.n288 w_19680_7310.n287 3.685
R3920 w_19680_7310.n282 w_19680_7310.n281 3.685
R3921 w_19680_7310.n276 w_19680_7310.n275 3.685
R3922 w_19680_7310.n270 w_19680_7310.n269 3.685
R3923 w_19680_7310.n48 w_19680_7310.n47 3.514
R3924 w_19680_7310.n264 w_19680_7310.n263 3.514
R3925 w_19680_7310.n399 w_19680_7310.n398 3.052
R3926 w_19680_7310.n393 w_19680_7310.n392 3.052
R3927 w_19680_7310.n387 w_19680_7310.n386 3.052
R3928 w_19680_7310.n381 w_19680_7310.n380 3.052
R3929 w_19680_7310.n375 w_19680_7310.n374 3.052
R3930 w_19680_7310.n370 w_19680_7310.n369 3.052
R3931 w_19680_7310.n363 w_19680_7310.n362 3.052
R3932 w_19680_7310.n357 w_19680_7310.n356 3.052
R3933 w_19680_7310.n351 w_19680_7310.n350 3.052
R3934 w_19680_7310.n345 w_19680_7310.n344 3.052
R3935 w_19680_7310.n475 w_19680_7310.n474 3.052
R3936 w_19680_7310.n469 w_19680_7310.n468 3.052
R3937 w_19680_7310.n463 w_19680_7310.n462 3.052
R3938 w_19680_7310.n457 w_19680_7310.n456 3.052
R3939 w_19680_7310.n451 w_19680_7310.n450 3.052
R3940 w_19680_7310.n446 w_19680_7310.n445 3.052
R3941 w_19680_7310.n439 w_19680_7310.n438 3.052
R3942 w_19680_7310.n433 w_19680_7310.n432 3.052
R3943 w_19680_7310.n427 w_19680_7310.n426 3.052
R3944 w_19680_7310.n421 w_19680_7310.n420 3.052
R3945 w_19680_7310.n510 w_19680_7310.n509 3.052
R3946 w_19680_7310.n516 w_19680_7310.n515 3.052
R3947 w_19680_7310.n522 w_19680_7310.n521 3.052
R3948 w_19680_7310.n528 w_19680_7310.n527 3.052
R3949 w_19680_7310.n37 w_19680_7310.n36 3.052
R3950 w_19680_7310.n2 w_19680_7310.n1 3.052
R3951 w_19680_7310.n30 w_19680_7310.n29 3.052
R3952 w_19680_7310.n24 w_19680_7310.n23 3.052
R3953 w_19680_7310.n18 w_19680_7310.n17 3.052
R3954 w_19680_7310.n12 w_19680_7310.n11 3.052
R3955 w_19680_7310.n178 w_19680_7310.n177 3.052
R3956 w_19680_7310.n172 w_19680_7310.n171 3.052
R3957 w_19680_7310.n166 w_19680_7310.n165 3.052
R3958 w_19680_7310.n160 w_19680_7310.n159 3.052
R3959 w_19680_7310.n154 w_19680_7310.n153 3.052
R3960 w_19680_7310.n149 w_19680_7310.n148 3.052
R3961 w_19680_7310.n142 w_19680_7310.n141 3.052
R3962 w_19680_7310.n136 w_19680_7310.n135 3.052
R3963 w_19680_7310.n130 w_19680_7310.n129 3.052
R3964 w_19680_7310.n124 w_19680_7310.n123 3.052
R3965 w_19680_7310.n339 w_19680_7310.n338 2.91
R3966 w_19680_7310.n415 w_19680_7310.n414 2.91
R3967 w_19680_7310.n6 w_19680_7310.n5 2.91
R3968 w_19680_7310.n118 w_19680_7310.n117 2.91
R3969 w_19680_7310.n189 w_19680_7310.n113 0.768
R3970 w_19680_7310.n410 w_19680_7310.n334 0.75
R3971 w_19680_7310.n52 w_19680_7310.n50 0.713
R3972 w_19680_7310.n196 w_19680_7310.n195 0.697
R3973 w_19680_7310.n196 w_19680_7310.n194 0.697
R3974 w_19680_7310.n197 w_19680_7310.n196 0.697
R3975 w_19680_7310.n196 w_19680_7310.n193 0.697
R3976 w_19680_7310.n196 w_19680_7310.n192 0.697
R3977 w_19680_7310.n196 w_19680_7310.n191 0.697
R3978 w_19680_7310.n268 w_19680_7310.n266 0.668
R3979 w_19680_7310.n205 w_19680_7310.n203 0.652
R3980 w_19680_7310.n10 w_19680_7310.n8 0.652
R3981 w_19680_7310.n343 w_19680_7310.n341 0.652
R3982 w_19680_7310.n419 w_19680_7310.n417 0.652
R3983 w_19680_7310.n122 w_19680_7310.n120 0.652
R3984 w_19680_7310.n42 w_19680_7310.n41 0.592
R3985 w_19680_7310.n486 w_19680_7310.n410 0.57
R3986 w_19680_7310.n259 w_19680_7310.n189 0.57
R3987 w_19680_7310.n498 w_19680_7310.n259 0.57
R3988 w_19680_7310.n498 w_19680_7310.n486 0.57
R3989 w_19680_7310.n410 w_19680_7310.n409 0.208
R3990 w_19680_7310.n486 w_19680_7310.n485 0.208
R3991 w_19680_7310.n189 w_19680_7310.n188 0.208
R3992 w_19680_7310.n259 w_19680_7310.n258 0.208
R3993 w_19680_7310.n501 w_19680_7310.n498 0.208
R3994 w_19680_7310.n489 w_19680_7310.n488 0.054
R3995 w_19680_7310.n491 w_19680_7310.n490 0.054
R3996 w_19680_7310.n493 w_19680_7310.n492 0.054
R3997 w_19680_7310.n495 w_19680_7310.n494 0.054
R3998 w_19680_7310.n497 w_19680_7310.n496 0.054
R3999 w_19680_7310.n304 w_19680_7310.n302 0.047
R4000 w_19680_7310.n80 w_19680_7310.n76 0.046
R4001 w_19680_7310.n113 w_19680_7310.n112 0.045
R4002 w_19680_7310.n488 w_19680_7310.n487 0.043
R4003 w_19680_7310.n490 w_19680_7310.n489 0.043
R4004 w_19680_7310.n492 w_19680_7310.n491 0.043
R4005 w_19680_7310.n494 w_19680_7310.n493 0.043
R4006 w_19680_7310.n496 w_19680_7310.n495 0.043
R4007 w_19680_7310.n297 w_19680_7310.n292 0.043
R4008 w_19680_7310.n84 w_19680_7310.n82 0.042
R4009 w_19680_7310.n334 w_19680_7310.n333 0.04
R4010 w_19680_7310.n333 w_19680_7310.n331 0.032
R4011 w_19680_7310.n331 w_19680_7310.n328 0.032
R4012 w_19680_7310.n328 w_19680_7310.n326 0.032
R4013 w_19680_7310.n326 w_19680_7310.n322 0.032
R4014 w_19680_7310.n322 w_19680_7310.n320 0.032
R4015 w_19680_7310.n320 w_19680_7310.n316 0.032
R4016 w_19680_7310.n316 w_19680_7310.n314 0.032
R4017 w_19680_7310.n314 w_19680_7310.n310 0.032
R4018 w_19680_7310.n310 w_19680_7310.n308 0.032
R4019 w_19680_7310.n308 w_19680_7310.n304 0.032
R4020 w_19680_7310.n292 w_19680_7310.n290 0.032
R4021 w_19680_7310.n290 w_19680_7310.n286 0.032
R4022 w_19680_7310.n286 w_19680_7310.n284 0.032
R4023 w_19680_7310.n284 w_19680_7310.n280 0.032
R4024 w_19680_7310.n280 w_19680_7310.n278 0.032
R4025 w_19680_7310.n278 w_19680_7310.n274 0.032
R4026 w_19680_7310.n274 w_19680_7310.n272 0.032
R4027 w_19680_7310.n272 w_19680_7310.n268 0.032
R4028 w_19680_7310.n379 w_19680_7310.n377 0.031
R4029 w_19680_7310.n455 w_19680_7310.n453 0.031
R4030 w_19680_7310.n158 w_19680_7310.n156 0.031
R4031 w_19680_7310.n232 w_19680_7310.n230 0.031
R4032 w_19680_7310.n533 w_19680_7310.n532 0.031
R4033 w_19680_7310.n112 w_19680_7310.n110 0.031
R4034 w_19680_7310.n110 w_19680_7310.n107 0.031
R4035 w_19680_7310.n107 w_19680_7310.n105 0.031
R4036 w_19680_7310.n105 w_19680_7310.n102 0.031
R4037 w_19680_7310.n102 w_19680_7310.n100 0.031
R4038 w_19680_7310.n100 w_19680_7310.n96 0.031
R4039 w_19680_7310.n96 w_19680_7310.n94 0.031
R4040 w_19680_7310.n94 w_19680_7310.n90 0.031
R4041 w_19680_7310.n90 w_19680_7310.n88 0.031
R4042 w_19680_7310.n88 w_19680_7310.n84 0.031
R4043 w_19680_7310.n76 w_19680_7310.n74 0.031
R4044 w_19680_7310.n74 w_19680_7310.n70 0.031
R4045 w_19680_7310.n70 w_19680_7310.n68 0.031
R4046 w_19680_7310.n68 w_19680_7310.n64 0.031
R4047 w_19680_7310.n64 w_19680_7310.n62 0.031
R4048 w_19680_7310.n62 w_19680_7310.n58 0.031
R4049 w_19680_7310.n58 w_19680_7310.n56 0.031
R4050 w_19680_7310.n56 w_19680_7310.n52 0.031
R4051 w_19680_7310.n302 w_19680_7310.n298 0.031
R4052 w_19680_7310.n81 w_19680_7310.n80 0.03
R4053 w_19680_7310.n372 w_19680_7310.n367 0.029
R4054 w_19680_7310.n448 w_19680_7310.n443 0.029
R4055 w_19680_7310.n151 w_19680_7310.n146 0.029
R4056 w_19680_7310.n226 w_19680_7310.n225 0.029
R4057 w_19680_7310.n35 w_19680_7310.n34 0.029
R4058 w_19680_7310.n409 w_19680_7310.n408 0.027
R4059 w_19680_7310.n485 w_19680_7310.n484 0.027
R4060 w_19680_7310.n188 w_19680_7310.n187 0.027
R4061 w_19680_7310.n258 w_19680_7310.n257 0.027
R4062 w_19680_7310.n503 w_19680_7310.n501 0.027
R4063 w_19680_7310.n408 w_19680_7310.n406 0.021
R4064 w_19680_7310.n406 w_19680_7310.n403 0.021
R4065 w_19680_7310.n403 w_19680_7310.n401 0.021
R4066 w_19680_7310.n401 w_19680_7310.n397 0.021
R4067 w_19680_7310.n397 w_19680_7310.n395 0.021
R4068 w_19680_7310.n395 w_19680_7310.n391 0.021
R4069 w_19680_7310.n391 w_19680_7310.n389 0.021
R4070 w_19680_7310.n389 w_19680_7310.n385 0.021
R4071 w_19680_7310.n385 w_19680_7310.n383 0.021
R4072 w_19680_7310.n383 w_19680_7310.n379 0.021
R4073 w_19680_7310.n367 w_19680_7310.n365 0.021
R4074 w_19680_7310.n365 w_19680_7310.n361 0.021
R4075 w_19680_7310.n361 w_19680_7310.n359 0.021
R4076 w_19680_7310.n359 w_19680_7310.n355 0.021
R4077 w_19680_7310.n355 w_19680_7310.n353 0.021
R4078 w_19680_7310.n353 w_19680_7310.n349 0.021
R4079 w_19680_7310.n349 w_19680_7310.n347 0.021
R4080 w_19680_7310.n347 w_19680_7310.n343 0.021
R4081 w_19680_7310.n484 w_19680_7310.n482 0.021
R4082 w_19680_7310.n482 w_19680_7310.n479 0.021
R4083 w_19680_7310.n479 w_19680_7310.n477 0.021
R4084 w_19680_7310.n477 w_19680_7310.n473 0.021
R4085 w_19680_7310.n473 w_19680_7310.n471 0.021
R4086 w_19680_7310.n471 w_19680_7310.n467 0.021
R4087 w_19680_7310.n467 w_19680_7310.n465 0.021
R4088 w_19680_7310.n465 w_19680_7310.n461 0.021
R4089 w_19680_7310.n461 w_19680_7310.n459 0.021
R4090 w_19680_7310.n459 w_19680_7310.n455 0.021
R4091 w_19680_7310.n443 w_19680_7310.n441 0.021
R4092 w_19680_7310.n441 w_19680_7310.n437 0.021
R4093 w_19680_7310.n437 w_19680_7310.n435 0.021
R4094 w_19680_7310.n435 w_19680_7310.n431 0.021
R4095 w_19680_7310.n431 w_19680_7310.n429 0.021
R4096 w_19680_7310.n429 w_19680_7310.n425 0.021
R4097 w_19680_7310.n425 w_19680_7310.n423 0.021
R4098 w_19680_7310.n423 w_19680_7310.n419 0.021
R4099 w_19680_7310.n187 w_19680_7310.n185 0.021
R4100 w_19680_7310.n185 w_19680_7310.n182 0.021
R4101 w_19680_7310.n182 w_19680_7310.n180 0.021
R4102 w_19680_7310.n180 w_19680_7310.n176 0.021
R4103 w_19680_7310.n176 w_19680_7310.n174 0.021
R4104 w_19680_7310.n174 w_19680_7310.n170 0.021
R4105 w_19680_7310.n170 w_19680_7310.n168 0.021
R4106 w_19680_7310.n168 w_19680_7310.n164 0.021
R4107 w_19680_7310.n164 w_19680_7310.n162 0.021
R4108 w_19680_7310.n162 w_19680_7310.n158 0.021
R4109 w_19680_7310.n146 w_19680_7310.n144 0.021
R4110 w_19680_7310.n144 w_19680_7310.n140 0.021
R4111 w_19680_7310.n140 w_19680_7310.n138 0.021
R4112 w_19680_7310.n138 w_19680_7310.n134 0.021
R4113 w_19680_7310.n134 w_19680_7310.n132 0.021
R4114 w_19680_7310.n132 w_19680_7310.n128 0.021
R4115 w_19680_7310.n128 w_19680_7310.n126 0.021
R4116 w_19680_7310.n126 w_19680_7310.n122 0.021
R4117 w_19680_7310.n257 w_19680_7310.n255 0.021
R4118 w_19680_7310.n255 w_19680_7310.n252 0.021
R4119 w_19680_7310.n252 w_19680_7310.n250 0.021
R4120 w_19680_7310.n250 w_19680_7310.n247 0.021
R4121 w_19680_7310.n247 w_19680_7310.n245 0.021
R4122 w_19680_7310.n245 w_19680_7310.n242 0.021
R4123 w_19680_7310.n242 w_19680_7310.n240 0.021
R4124 w_19680_7310.n240 w_19680_7310.n237 0.021
R4125 w_19680_7310.n237 w_19680_7310.n235 0.021
R4126 w_19680_7310.n235 w_19680_7310.n232 0.021
R4127 w_19680_7310.n225 w_19680_7310.n223 0.021
R4128 w_19680_7310.n223 w_19680_7310.n220 0.021
R4129 w_19680_7310.n220 w_19680_7310.n218 0.021
R4130 w_19680_7310.n218 w_19680_7310.n215 0.021
R4131 w_19680_7310.n215 w_19680_7310.n213 0.021
R4132 w_19680_7310.n213 w_19680_7310.n210 0.021
R4133 w_19680_7310.n210 w_19680_7310.n208 0.021
R4134 w_19680_7310.n208 w_19680_7310.n205 0.021
R4135 w_19680_7310.n506 w_19680_7310.n503 0.021
R4136 w_19680_7310.n508 w_19680_7310.n506 0.021
R4137 w_19680_7310.n512 w_19680_7310.n508 0.021
R4138 w_19680_7310.n514 w_19680_7310.n512 0.021
R4139 w_19680_7310.n518 w_19680_7310.n514 0.021
R4140 w_19680_7310.n520 w_19680_7310.n518 0.021
R4141 w_19680_7310.n524 w_19680_7310.n520 0.021
R4142 w_19680_7310.n526 w_19680_7310.n524 0.021
R4143 w_19680_7310.n530 w_19680_7310.n526 0.021
R4144 w_19680_7310.n532 w_19680_7310.n530 0.021
R4145 w_19680_7310.n34 w_19680_7310.n32 0.021
R4146 w_19680_7310.n32 w_19680_7310.n28 0.021
R4147 w_19680_7310.n28 w_19680_7310.n26 0.021
R4148 w_19680_7310.n26 w_19680_7310.n22 0.021
R4149 w_19680_7310.n22 w_19680_7310.n20 0.021
R4150 w_19680_7310.n20 w_19680_7310.n16 0.021
R4151 w_19680_7310.n16 w_19680_7310.n14 0.021
R4152 w_19680_7310.n14 w_19680_7310.n10 0.021
R4153 w_19680_7310.n377 w_19680_7310.n373 0.021
R4154 w_19680_7310.n453 w_19680_7310.n449 0.021
R4155 w_19680_7310.n534 w_19680_7310.n533 0.021
R4156 w_19680_7310.n156 w_19680_7310.n152 0.021
R4157 w_19680_7310.n230 w_19680_7310.n227 0.021
R4158 w_19680_7310.n298 w_19680_7310.n297 0.009
R4159 w_19680_7310.n82 w_19680_7310.n81 0.009
R4160 w_19680_7310.n373 w_19680_7310.n372 0.006
R4161 w_19680_7310.n449 w_19680_7310.n448 0.006
R4162 w_19680_7310.n534 w_19680_7310.n35 0.006
R4163 w_19680_7310.n152 w_19680_7310.n151 0.006
R4164 w_19680_7310.n227 w_19680_7310.n226 0.006
C0 vrec vinn 0.80fF
C1 vrec vinp 1.14fF
C2 vinn vinp 14.67fF
.ends

