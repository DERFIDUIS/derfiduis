magic
tech sky130A
magscale 1 2
timestamp 1680449562
<< xpolycontact >>
rect -35 1410 35 1842
rect -35 -1842 35 -1410
<< xpolyres >>
rect -35 -1410 35 1410
<< viali >>
rect -19 1427 19 1824
rect -19 -1824 19 -1427
<< metal1 >>
rect -25 1824 25 1836
rect -25 1427 -19 1824
rect 19 1427 25 1824
rect -25 1415 25 1427
rect -25 -1427 25 -1415
rect -25 -1824 -19 -1427
rect 19 -1824 25 -1427
rect -25 -1836 25 -1824
<< res1p41 >>
rect -37 -1412 37 1412
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 0.350 l 14.1 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 81.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
