magic
tech sky130A
timestamp 1680257378
<< pwell >>
rect -448 -355 448 355
<< nmoslvt >>
rect -350 -250 350 250
<< ndiff >>
rect -379 244 -350 250
rect -379 -244 -373 244
rect -356 -244 -350 244
rect -379 -250 -350 -244
rect 350 244 379 250
rect 350 -244 356 244
rect 373 -244 379 244
rect 350 -250 379 -244
<< ndiffc >>
rect -373 -244 -356 244
rect 356 -244 373 244
<< psubdiff >>
rect -430 320 -382 337
rect 382 320 430 337
rect -430 289 -413 320
rect 413 289 430 320
rect -430 -320 -413 -289
rect 413 -320 430 -289
rect -430 -337 -382 -320
rect 382 -337 430 -320
<< psubdiffcont >>
rect -382 320 382 337
rect -430 -289 -413 289
rect 413 -289 430 289
rect -382 -337 382 -320
<< poly >>
rect -350 286 350 294
rect -350 269 -342 286
rect 342 269 350 286
rect -350 250 350 269
rect -350 -269 350 -250
rect -350 -286 -342 -269
rect 342 -286 350 -269
rect -350 -294 350 -286
<< polycont >>
rect -342 269 342 286
rect -342 -286 342 -269
<< locali >>
rect -430 320 -382 337
rect 382 320 430 337
rect -430 289 -413 320
rect 413 289 430 320
rect -350 269 -342 286
rect 342 269 350 286
rect -373 244 -356 252
rect -373 -252 -356 -244
rect 356 244 373 252
rect 356 -252 373 -244
rect -350 -286 -342 -269
rect 342 -286 350 -269
rect -430 -320 -413 -289
rect 413 -320 430 -289
rect -430 -337 -382 -320
rect 382 -337 430 -320
<< viali >>
rect -342 269 342 286
rect -373 -244 -356 244
rect 356 -244 373 244
rect -342 -286 342 -269
<< metal1 >>
rect -348 286 348 289
rect -348 269 -342 286
rect 342 269 348 286
rect -348 266 348 269
rect -376 244 -353 250
rect -376 -244 -373 244
rect -356 -244 -353 244
rect -376 -250 -353 -244
rect 353 244 376 250
rect 353 -244 356 244
rect 373 -244 376 244
rect 353 -250 376 -244
rect -348 -269 348 -266
rect -348 -286 -342 -269
rect 342 -286 348 -269
rect -348 -289 348 -286
<< properties >>
string FIXED_BBOX -421 -328 421 328
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.0 l 7.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
