magic
tech sky130A
magscale 1 2
timestamp 1681673980
<< nwell >>
rect -294 -864 294 898
<< pmoslvt >>
rect -200 -764 200 836
<< pdiff >>
rect -258 824 -200 836
rect -258 -752 -246 824
rect -212 -752 -200 824
rect -258 -764 -200 -752
rect 200 824 258 836
rect 200 -752 212 824
rect 246 -752 258 824
rect 200 -764 258 -752
<< pdiffc >>
rect -246 -752 -212 824
rect 212 -752 246 824
<< poly >>
rect -200 836 200 862
rect -200 -811 200 -764
rect -200 -845 -184 -811
rect 184 -845 200 -811
rect -200 -861 200 -845
<< polycont >>
rect -184 -845 184 -811
<< locali >>
rect -246 824 -212 840
rect -246 -768 -212 -752
rect 212 824 246 840
rect 212 -768 246 -752
rect -200 -845 -184 -811
rect 184 -845 200 -811
<< viali >>
rect -246 -752 -212 824
rect 212 -752 246 824
rect -184 -845 184 -811
<< metal1 >>
rect -252 824 -206 836
rect -252 -752 -246 824
rect -212 -752 -206 824
rect -252 -764 -206 -752
rect 206 824 252 836
rect 206 -752 212 824
rect 246 -752 252 824
rect 206 -764 252 -752
rect -196 -811 196 -805
rect -196 -845 -184 -811
rect 184 -845 196 -811
rect -196 -851 196 -845
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 8.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
