magic
tech sky130A
magscale 1 2
timestamp 1682034855
<< metal4 >>
rect -2909 2599 2909 2640
rect -2909 -2599 2653 2599
rect 2889 -2599 2909 2599
rect -2909 -2640 2909 -2599
<< via4 >>
rect 2653 -2599 2889 2599
<< mimcap2 >>
rect -2829 2520 2291 2560
rect -2829 -2520 -2789 2520
rect 2251 -2520 2291 2520
rect -2829 -2560 2291 -2520
<< mimcap2contact >>
rect -2789 -2520 2251 2520
<< metal5 >>
rect 2611 2599 2931 2641
rect -2813 2520 2275 2544
rect -2813 -2520 -2789 2520
rect 2251 -2520 2275 2520
rect -2813 -2544 2275 -2520
rect 2611 -2599 2653 2599
rect 2889 -2599 2931 2599
rect 2611 -2641 2931 -2599
<< properties >>
string FIXED_BBOX -2909 -2640 2371 2640
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25.6 l 25.6 val 1.33k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
