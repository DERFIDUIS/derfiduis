* NGSPICE file created from Temperature_Sensor.ext - technology: sky130A

.subckt Temperature_Sensor vtemp iin vdd vss
M61 a_n3070_n3662# a_n4954_n2108# vdd vss sky130_fd_pr__nfet_01v8_lvt ad=1.2e+13p pd=8.6e+07u as=1.843e+13p ps=1.1424e+08u w=4e+06u l=2e+06u
M71 a_62_n3936# a_n3216_n2108# a_n178_n2405# vss sky130_fd_pr__nfet_01v8_lvt ad=1.635e+13p pd=1.1654e+08u as=2.9e+12p ps=2.116e+07u w=5e+06u l=2e+06u
M62 a_n3070_n3662# a_n4954_n2108# vdd vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
M94 a_n178_n2405# a_n178_n2405# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=2.9e+12p pd=2.116e+07u as=1.44e+13p ps=1.02e+08u w=5e+06u l=2e+06u
M2 a_n4896_n2205# iin vss vss sky130_fd_pr__nfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=1.33825e+13p ps=8.728e+07u w=4e+06u l=2e+06u
M81 vtemp a_n3070_n3662# a_62_n3936# vss sky130_fd_pr__nfet_01v8_lvt ad=2.9e+12p pd=2.116e+07u as=0p ps=0u w=5e+06u l=500000u
M72 a_n178_n2405# a_n3216_n2108# a_62_n3936# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M73 a_n178_n2405# a_n3216_n2108# a_62_n3936# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M5 a_n3216_n2108# a_n4954_n2108# a_n4954_n2108# vss sky130_fd_pr__nfet_01v8_lvt ad=1.2e+12p pd=8.6e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=2e+06u
M93 vdd a_n178_n2405# a_n178_n2405# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M63 vdd a_n4954_n2108# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
M82 a_62_n3936# a_n3070_n3662# vtemp vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
M92 a_n178_n2405# a_n178_n2405# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M64 vdd a_n4954_n2108# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
M65 vdd a_n4954_n2108# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
M83 a_62_n3936# a_n3070_n3662# vtemp vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
M112 vss iin a_62_n3936# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M111 vss iin a_62_n3936# vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M66 a_n3070_n3662# a_n4954_n2108# vdd vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
Q3 vss vss a_n3216_n2108# sky130_fd_pr__pnp_05v5_W3p40L3p40
M3 a_n4896_n2205# a_n4896_n2205# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=1.16e+12p pd=8.58e+06u as=0p ps=0u w=4e+06u l=2e+06u
M1 vss iin iin vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=2e+06u
M104 vdd a_n178_n2405# vtemp vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+12p ps=2.116e+07u w=5e+06u l=2e+06u
M103 vtemp a_n178_n2405# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M67 a_n3070_n3662# a_n4954_n2108# vdd vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
Q4 vss vss a_n3070_n3662# sky130_fd_pr__pnp_05v5_W3p40L3p40
M113 a_62_n3936# iin vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M68 vdd a_n4954_n2108# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
M69 vdd a_n4954_n2108# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
M84 vtemp a_n3070_n3662# a_62_n3936# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
M74 a_62_n3936# a_n3216_n2108# a_n178_n2405# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M102 vtemp a_n178_n2405# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M101 vdd a_n178_n2405# vtemp vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M4 vdd a_n4896_n2205# a_n4954_n2108# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.16e+12p ps=8.58e+06u w=4e+06u l=2e+06u
M91 vdd a_n178_n2405# a_n178_n2405# vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
M610 vdd a_n4954_n2108# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
M114 a_62_n3936# iin vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
.ends

