magic
tech sky130A
magscale 1 2
timestamp 1681578886
<< nwell >>
rect -4902 -2072 -4898 -2064
rect -4450 -2208 -4336 -1246
rect -3906 -2198 -3890 -2146
rect -340 -2302 -224 -1246
rect -340 -2408 -174 -2302
rect 726 -2408 840 -1246
rect 1790 -2408 1904 -1246
rect 2854 -2408 2968 -1246
rect 3930 -2408 4034 -1246
<< nbase >>
rect -2770 -4356 -2742 -4316
rect -2480 -4322 -2466 -4316
rect -2486 -4356 -2466 -4322
rect -1630 -4332 -1622 -4296
rect -1574 -4356 -1556 -4322
rect -2766 -4392 -2762 -4356
rect -2770 -4524 -2726 -4392
rect -2766 -4532 -2762 -4524
rect -2766 -4600 -2760 -4532
rect -2480 -4600 -2472 -4356
rect -1572 -4392 -1568 -4356
rect -1578 -4524 -1558 -4392
rect -1572 -4592 -1568 -4524
rect -1572 -4600 -1566 -4592
rect -1290 -4600 -1284 -4592
rect -2766 -4606 -2474 -4600
rect -1572 -4606 -1284 -4600
<< ndiff >>
rect -3158 -2108 -3156 -1308
rect -3070 -2108 -3068 -1308
rect -2094 -2108 -2092 -1308
rect -2006 -2108 -2004 -1308
rect -1030 -2108 -1028 -1308
rect -942 -2108 -940 -1308
rect -4438 -3662 -4436 -2862
rect -4350 -3662 -4348 -2862
rect -3070 -3662 -3068 -2862
rect -2094 -3662 -2092 -2862
rect -2006 -3662 -2004 -2862
rect -1030 -3662 -1028 -2862
rect -942 -3662 -940 -2862
rect 62 -3936 64 -2936
rect 438 -3936 440 -2936
rect 526 -3936 528 -2936
rect 1502 -3936 1504 -2936
rect 2190 -3936 2192 -2936
rect 2566 -3936 2568 -2936
rect 2654 -3936 2656 -2936
rect 3630 -3936 3632 -2936
rect 1264 -5384 1266 -4384
rect 1352 -5384 1354 -4384
rect 2328 -5384 2330 -4384
rect 2416 -5384 2418 -4384
<< pdiff >>
rect -4902 -2072 -4898 -2064
rect -4438 -2108 -4436 -1308
rect -4350 -2108 -4348 -1308
rect -238 -2308 -236 -1308
rect 738 -2308 740 -1308
rect 826 -2308 828 -1308
rect 1802 -2308 1804 -1308
rect 1890 -2308 1892 -1308
rect 2866 -2308 2868 -1308
rect 2954 -2308 2956 -1308
rect 3930 -2308 3932 -1308
<< psubdiff >>
rect -3156 -1366 -3070 -1308
rect -3156 -1400 -3130 -1366
rect -3096 -1400 -3070 -1366
rect -3156 -1434 -3070 -1400
rect -3156 -1468 -3130 -1434
rect -3096 -1468 -3070 -1434
rect -3156 -1502 -3070 -1468
rect -3156 -1536 -3130 -1502
rect -3096 -1536 -3070 -1502
rect -3156 -1570 -3070 -1536
rect -3156 -1604 -3130 -1570
rect -3096 -1604 -3070 -1570
rect -3156 -1638 -3070 -1604
rect -3156 -1672 -3130 -1638
rect -3096 -1672 -3070 -1638
rect -3156 -1706 -3070 -1672
rect -3156 -1740 -3130 -1706
rect -3096 -1740 -3070 -1706
rect -3156 -1774 -3070 -1740
rect -3156 -1808 -3130 -1774
rect -3096 -1808 -3070 -1774
rect -3156 -1842 -3070 -1808
rect -3156 -1876 -3130 -1842
rect -3096 -1876 -3070 -1842
rect -3156 -1910 -3070 -1876
rect -3156 -1944 -3130 -1910
rect -3096 -1944 -3070 -1910
rect -3156 -1978 -3070 -1944
rect -3156 -2012 -3130 -1978
rect -3096 -2012 -3070 -1978
rect -3156 -2046 -3070 -2012
rect -3156 -2080 -3130 -2046
rect -3096 -2080 -3070 -2046
rect -3156 -2108 -3070 -2080
rect -2092 -1366 -2006 -1308
rect -2092 -1400 -2066 -1366
rect -2032 -1400 -2006 -1366
rect -2092 -1434 -2006 -1400
rect -2092 -1468 -2066 -1434
rect -2032 -1468 -2006 -1434
rect -2092 -1502 -2006 -1468
rect -2092 -1536 -2066 -1502
rect -2032 -1536 -2006 -1502
rect -2092 -1570 -2006 -1536
rect -2092 -1604 -2066 -1570
rect -2032 -1604 -2006 -1570
rect -2092 -1638 -2006 -1604
rect -2092 -1672 -2066 -1638
rect -2032 -1672 -2006 -1638
rect -2092 -1706 -2006 -1672
rect -2092 -1740 -2066 -1706
rect -2032 -1740 -2006 -1706
rect -2092 -1774 -2006 -1740
rect -2092 -1808 -2066 -1774
rect -2032 -1808 -2006 -1774
rect -2092 -1842 -2006 -1808
rect -2092 -1876 -2066 -1842
rect -2032 -1876 -2006 -1842
rect -2092 -1910 -2006 -1876
rect -2092 -1944 -2066 -1910
rect -2032 -1944 -2006 -1910
rect -2092 -1978 -2006 -1944
rect -2092 -2012 -2066 -1978
rect -2032 -2012 -2006 -1978
rect -2092 -2046 -2006 -2012
rect -2092 -2080 -2066 -2046
rect -2032 -2080 -2006 -2046
rect -2092 -2108 -2006 -2080
rect -1028 -1366 -942 -1308
rect -1028 -1400 -1002 -1366
rect -968 -1400 -942 -1366
rect -1028 -1434 -942 -1400
rect -1028 -1468 -1002 -1434
rect -968 -1468 -942 -1434
rect -1028 -1502 -942 -1468
rect -1028 -1536 -1002 -1502
rect -968 -1536 -942 -1502
rect -1028 -1570 -942 -1536
rect -1028 -1604 -1002 -1570
rect -968 -1604 -942 -1570
rect -1028 -1638 -942 -1604
rect -1028 -1672 -1002 -1638
rect -968 -1672 -942 -1638
rect -1028 -1706 -942 -1672
rect -1028 -1740 -1002 -1706
rect -968 -1740 -942 -1706
rect -1028 -1774 -942 -1740
rect -1028 -1808 -1002 -1774
rect -968 -1808 -942 -1774
rect -1028 -1842 -942 -1808
rect -1028 -1876 -1002 -1842
rect -968 -1876 -942 -1842
rect -1028 -1910 -942 -1876
rect -1028 -1944 -1002 -1910
rect -968 -1944 -942 -1910
rect -1028 -1978 -942 -1944
rect -1028 -2012 -1002 -1978
rect -968 -2012 -942 -1978
rect -1028 -2046 -942 -2012
rect -1028 -2080 -1002 -2046
rect -968 -2080 -942 -2046
rect -1028 -2108 -942 -2080
rect -4436 -2920 -4350 -2862
rect -4436 -2954 -4410 -2920
rect -4376 -2954 -4350 -2920
rect -4436 -2988 -4350 -2954
rect -4436 -3022 -4410 -2988
rect -4376 -3022 -4350 -2988
rect -4436 -3056 -4350 -3022
rect -4436 -3090 -4410 -3056
rect -4376 -3090 -4350 -3056
rect -4436 -3124 -4350 -3090
rect -4436 -3158 -4410 -3124
rect -4376 -3158 -4350 -3124
rect -4436 -3192 -4350 -3158
rect -4436 -3226 -4410 -3192
rect -4376 -3226 -4350 -3192
rect -4436 -3260 -4350 -3226
rect -4436 -3294 -4410 -3260
rect -4376 -3294 -4350 -3260
rect -4436 -3328 -4350 -3294
rect -4436 -3362 -4410 -3328
rect -4376 -3362 -4350 -3328
rect -4436 -3396 -4350 -3362
rect -4436 -3430 -4410 -3396
rect -4376 -3430 -4350 -3396
rect -4436 -3464 -4350 -3430
rect -4436 -3498 -4410 -3464
rect -4376 -3498 -4350 -3464
rect -4436 -3532 -4350 -3498
rect -4436 -3566 -4410 -3532
rect -4376 -3566 -4350 -3532
rect -4436 -3600 -4350 -3566
rect -4436 -3634 -4410 -3600
rect -4376 -3634 -4350 -3600
rect -4436 -3662 -4350 -3634
rect -3134 -2920 -3070 -2862
rect -3134 -2954 -3130 -2920
rect -3096 -2954 -3070 -2920
rect -3134 -2988 -3070 -2954
rect -3134 -3022 -3130 -2988
rect -3096 -3022 -3070 -2988
rect -3134 -3056 -3070 -3022
rect -3134 -3090 -3130 -3056
rect -3096 -3090 -3070 -3056
rect -3134 -3124 -3070 -3090
rect -3134 -3158 -3130 -3124
rect -3096 -3158 -3070 -3124
rect -3134 -3192 -3070 -3158
rect -3134 -3226 -3130 -3192
rect -3096 -3226 -3070 -3192
rect -3134 -3260 -3070 -3226
rect -3134 -3294 -3130 -3260
rect -3096 -3294 -3070 -3260
rect -3134 -3328 -3070 -3294
rect -3134 -3362 -3130 -3328
rect -3096 -3362 -3070 -3328
rect -3134 -3396 -3070 -3362
rect -3134 -3430 -3130 -3396
rect -3096 -3430 -3070 -3396
rect -3134 -3464 -3070 -3430
rect -3134 -3498 -3130 -3464
rect -3096 -3498 -3070 -3464
rect -3134 -3532 -3070 -3498
rect -3134 -3566 -3130 -3532
rect -3096 -3566 -3070 -3532
rect -3134 -3600 -3070 -3566
rect -3134 -3634 -3130 -3600
rect -3096 -3634 -3070 -3600
rect -3134 -3662 -3070 -3634
rect -2092 -2920 -2006 -2862
rect -2092 -2954 -2066 -2920
rect -2032 -2954 -2006 -2920
rect -2092 -2988 -2006 -2954
rect -2092 -3022 -2066 -2988
rect -2032 -3022 -2006 -2988
rect -2092 -3056 -2006 -3022
rect -2092 -3090 -2066 -3056
rect -2032 -3090 -2006 -3056
rect -2092 -3124 -2006 -3090
rect -2092 -3158 -2066 -3124
rect -2032 -3158 -2006 -3124
rect -2092 -3192 -2006 -3158
rect -2092 -3226 -2066 -3192
rect -2032 -3226 -2006 -3192
rect -2092 -3260 -2006 -3226
rect -2092 -3294 -2066 -3260
rect -2032 -3294 -2006 -3260
rect -2092 -3328 -2006 -3294
rect -2092 -3362 -2066 -3328
rect -2032 -3362 -2006 -3328
rect -2092 -3396 -2006 -3362
rect -2092 -3430 -2066 -3396
rect -2032 -3430 -2006 -3396
rect -2092 -3464 -2006 -3430
rect -2092 -3498 -2066 -3464
rect -2032 -3498 -2006 -3464
rect -2092 -3532 -2006 -3498
rect -2092 -3566 -2066 -3532
rect -2032 -3566 -2006 -3532
rect -2092 -3600 -2006 -3566
rect -2092 -3634 -2066 -3600
rect -2032 -3634 -2006 -3600
rect -2092 -3662 -2006 -3634
rect -1028 -2920 -942 -2862
rect -1028 -2954 -1002 -2920
rect -968 -2954 -942 -2920
rect -1028 -2988 -942 -2954
rect -1028 -3022 -1002 -2988
rect -968 -3022 -942 -2988
rect -1028 -3056 -942 -3022
rect -1028 -3090 -1002 -3056
rect -968 -3090 -942 -3056
rect -1028 -3124 -942 -3090
rect -1028 -3158 -1002 -3124
rect -968 -3158 -942 -3124
rect -1028 -3192 -942 -3158
rect -1028 -3226 -1002 -3192
rect -968 -3226 -942 -3192
rect -1028 -3260 -942 -3226
rect -1028 -3294 -1002 -3260
rect -968 -3294 -942 -3260
rect -1028 -3328 -942 -3294
rect -1028 -3362 -1002 -3328
rect -968 -3362 -942 -3328
rect -1028 -3396 -942 -3362
rect -1028 -3430 -1002 -3396
rect -968 -3430 -942 -3396
rect -1028 -3464 -942 -3430
rect -1028 -3498 -1002 -3464
rect -968 -3498 -942 -3464
rect -1028 -3532 -942 -3498
rect -1028 -3566 -1002 -3532
rect -968 -3566 -942 -3532
rect -1028 -3600 -942 -3566
rect -1028 -3634 -1002 -3600
rect -968 -3634 -942 -3600
rect -1028 -3662 -942 -3634
rect -2 -2990 62 -2936
rect -2 -3024 2 -2990
rect 36 -3024 62 -2990
rect -2 -3058 62 -3024
rect -2 -3092 2 -3058
rect 36 -3092 62 -3058
rect -2 -3126 62 -3092
rect -2 -3160 2 -3126
rect 36 -3160 62 -3126
rect -2 -3194 62 -3160
rect -2 -3228 2 -3194
rect 36 -3228 62 -3194
rect -2 -3262 62 -3228
rect -2 -3296 2 -3262
rect 36 -3296 62 -3262
rect -2 -3330 62 -3296
rect -2 -3364 2 -3330
rect 36 -3364 62 -3330
rect -2 -3398 62 -3364
rect -2 -3432 2 -3398
rect 36 -3432 62 -3398
rect -2 -3466 62 -3432
rect -2 -3500 2 -3466
rect 36 -3500 62 -3466
rect -2 -3534 62 -3500
rect -2 -3568 2 -3534
rect 36 -3568 62 -3534
rect -2 -3602 62 -3568
rect -2 -3636 2 -3602
rect 36 -3636 62 -3602
rect -2 -3670 62 -3636
rect -2 -3704 2 -3670
rect 36 -3704 62 -3670
rect -2 -3738 62 -3704
rect -2 -3772 2 -3738
rect 36 -3772 62 -3738
rect -2 -3806 62 -3772
rect -2 -3840 2 -3806
rect 36 -3840 62 -3806
rect -2 -3874 62 -3840
rect -2 -3908 2 -3874
rect 36 -3908 62 -3874
rect -2 -3936 62 -3908
rect 440 -2990 526 -2936
rect 440 -3024 466 -2990
rect 500 -3024 526 -2990
rect 440 -3058 526 -3024
rect 440 -3092 466 -3058
rect 500 -3092 526 -3058
rect 440 -3126 526 -3092
rect 440 -3160 466 -3126
rect 500 -3160 526 -3126
rect 440 -3194 526 -3160
rect 440 -3228 466 -3194
rect 500 -3228 526 -3194
rect 440 -3262 526 -3228
rect 440 -3296 466 -3262
rect 500 -3296 526 -3262
rect 440 -3330 526 -3296
rect 440 -3364 466 -3330
rect 500 -3364 526 -3330
rect 440 -3398 526 -3364
rect 440 -3432 466 -3398
rect 500 -3432 526 -3398
rect 440 -3466 526 -3432
rect 440 -3500 466 -3466
rect 500 -3500 526 -3466
rect 440 -3534 526 -3500
rect 440 -3568 466 -3534
rect 500 -3568 526 -3534
rect 440 -3602 526 -3568
rect 440 -3636 466 -3602
rect 500 -3636 526 -3602
rect 440 -3670 526 -3636
rect 440 -3704 466 -3670
rect 500 -3704 526 -3670
rect 440 -3738 526 -3704
rect 440 -3772 466 -3738
rect 500 -3772 526 -3738
rect 440 -3806 526 -3772
rect 440 -3840 466 -3806
rect 500 -3840 526 -3806
rect 440 -3874 526 -3840
rect 440 -3908 466 -3874
rect 500 -3908 526 -3874
rect 440 -3936 526 -3908
rect 1504 -2990 1570 -2936
rect 1504 -3024 1530 -2990
rect 1564 -3024 1570 -2990
rect 1504 -3058 1570 -3024
rect 1504 -3092 1530 -3058
rect 1564 -3092 1570 -3058
rect 1504 -3126 1570 -3092
rect 1504 -3160 1530 -3126
rect 1564 -3160 1570 -3126
rect 1504 -3194 1570 -3160
rect 1504 -3228 1530 -3194
rect 1564 -3228 1570 -3194
rect 1504 -3262 1570 -3228
rect 1504 -3296 1530 -3262
rect 1564 -3296 1570 -3262
rect 1504 -3330 1570 -3296
rect 1504 -3364 1530 -3330
rect 1564 -3364 1570 -3330
rect 1504 -3398 1570 -3364
rect 1504 -3432 1530 -3398
rect 1564 -3432 1570 -3398
rect 1504 -3466 1570 -3432
rect 1504 -3500 1530 -3466
rect 1564 -3500 1570 -3466
rect 1504 -3534 1570 -3500
rect 1504 -3568 1530 -3534
rect 1564 -3568 1570 -3534
rect 1504 -3602 1570 -3568
rect 1504 -3636 1530 -3602
rect 1564 -3636 1570 -3602
rect 1504 -3670 1570 -3636
rect 1504 -3704 1530 -3670
rect 1564 -3704 1570 -3670
rect 1504 -3738 1570 -3704
rect 1504 -3772 1530 -3738
rect 1564 -3772 1570 -3738
rect 1504 -3806 1570 -3772
rect 1504 -3840 1530 -3806
rect 1564 -3840 1570 -3806
rect 1504 -3874 1570 -3840
rect 1504 -3908 1530 -3874
rect 1564 -3908 1570 -3874
rect 1504 -3936 1570 -3908
rect 2124 -2990 2190 -2936
rect 2124 -3024 2130 -2990
rect 2164 -3024 2190 -2990
rect 2124 -3058 2190 -3024
rect 2124 -3092 2130 -3058
rect 2164 -3092 2190 -3058
rect 2124 -3126 2190 -3092
rect 2124 -3160 2130 -3126
rect 2164 -3160 2190 -3126
rect 2124 -3194 2190 -3160
rect 2124 -3228 2130 -3194
rect 2164 -3228 2190 -3194
rect 2124 -3262 2190 -3228
rect 2124 -3296 2130 -3262
rect 2164 -3296 2190 -3262
rect 2124 -3330 2190 -3296
rect 2124 -3364 2130 -3330
rect 2164 -3364 2190 -3330
rect 2124 -3398 2190 -3364
rect 2124 -3432 2130 -3398
rect 2164 -3432 2190 -3398
rect 2124 -3466 2190 -3432
rect 2124 -3500 2130 -3466
rect 2164 -3500 2190 -3466
rect 2124 -3534 2190 -3500
rect 2124 -3568 2130 -3534
rect 2164 -3568 2190 -3534
rect 2124 -3602 2190 -3568
rect 2124 -3636 2130 -3602
rect 2164 -3636 2190 -3602
rect 2124 -3670 2190 -3636
rect 2124 -3704 2130 -3670
rect 2164 -3704 2190 -3670
rect 2124 -3738 2190 -3704
rect 2124 -3772 2130 -3738
rect 2164 -3772 2190 -3738
rect 2124 -3806 2190 -3772
rect 2124 -3840 2130 -3806
rect 2164 -3840 2190 -3806
rect 2124 -3874 2190 -3840
rect 2124 -3908 2130 -3874
rect 2164 -3908 2190 -3874
rect 2124 -3936 2190 -3908
rect 2568 -2990 2654 -2936
rect 2568 -3024 2594 -2990
rect 2628 -3024 2654 -2990
rect 2568 -3058 2654 -3024
rect 2568 -3092 2594 -3058
rect 2628 -3092 2654 -3058
rect 2568 -3126 2654 -3092
rect 2568 -3160 2594 -3126
rect 2628 -3160 2654 -3126
rect 2568 -3194 2654 -3160
rect 2568 -3228 2594 -3194
rect 2628 -3228 2654 -3194
rect 2568 -3262 2654 -3228
rect 2568 -3296 2594 -3262
rect 2628 -3296 2654 -3262
rect 2568 -3330 2654 -3296
rect 2568 -3364 2594 -3330
rect 2628 -3364 2654 -3330
rect 2568 -3398 2654 -3364
rect 2568 -3432 2594 -3398
rect 2628 -3432 2654 -3398
rect 2568 -3466 2654 -3432
rect 2568 -3500 2594 -3466
rect 2628 -3500 2654 -3466
rect 2568 -3534 2654 -3500
rect 2568 -3568 2594 -3534
rect 2628 -3568 2654 -3534
rect 2568 -3602 2654 -3568
rect 2568 -3636 2594 -3602
rect 2628 -3636 2654 -3602
rect 2568 -3670 2654 -3636
rect 2568 -3704 2594 -3670
rect 2628 -3704 2654 -3670
rect 2568 -3738 2654 -3704
rect 2568 -3772 2594 -3738
rect 2628 -3772 2654 -3738
rect 2568 -3806 2654 -3772
rect 2568 -3840 2594 -3806
rect 2628 -3840 2654 -3806
rect 2568 -3874 2654 -3840
rect 2568 -3908 2594 -3874
rect 2628 -3908 2654 -3874
rect 2568 -3936 2654 -3908
rect 3632 -2990 3696 -2936
rect 3632 -3024 3658 -2990
rect 3692 -3024 3696 -2990
rect 3632 -3058 3696 -3024
rect 3632 -3092 3658 -3058
rect 3692 -3092 3696 -3058
rect 3632 -3126 3696 -3092
rect 3632 -3160 3658 -3126
rect 3692 -3160 3696 -3126
rect 3632 -3194 3696 -3160
rect 3632 -3228 3658 -3194
rect 3692 -3228 3696 -3194
rect 3632 -3262 3696 -3228
rect 3632 -3296 3658 -3262
rect 3692 -3296 3696 -3262
rect 3632 -3330 3696 -3296
rect 3632 -3364 3658 -3330
rect 3692 -3364 3696 -3330
rect 3632 -3398 3696 -3364
rect 3632 -3432 3658 -3398
rect 3692 -3432 3696 -3398
rect 3632 -3466 3696 -3432
rect 3632 -3500 3658 -3466
rect 3692 -3500 3696 -3466
rect 3632 -3534 3696 -3500
rect 3632 -3568 3658 -3534
rect 3692 -3568 3696 -3534
rect 3632 -3602 3696 -3568
rect 3632 -3636 3658 -3602
rect 3692 -3636 3696 -3602
rect 3632 -3670 3696 -3636
rect 3632 -3704 3658 -3670
rect 3692 -3704 3696 -3670
rect 3632 -3738 3696 -3704
rect 3632 -3772 3658 -3738
rect 3692 -3772 3696 -3738
rect 3632 -3806 3696 -3772
rect 3632 -3840 3658 -3806
rect 3692 -3840 3696 -3806
rect 3632 -3874 3696 -3840
rect 3632 -3908 3658 -3874
rect 3692 -3908 3696 -3874
rect 3632 -3936 3696 -3908
rect 1266 -4438 1352 -4384
rect 1266 -4472 1292 -4438
rect 1326 -4472 1352 -4438
rect 1266 -4506 1352 -4472
rect 1266 -4540 1292 -4506
rect 1326 -4540 1352 -4506
rect 1266 -4574 1352 -4540
rect 1266 -4608 1292 -4574
rect 1326 -4608 1352 -4574
rect 1266 -4642 1352 -4608
rect 1266 -4676 1292 -4642
rect 1326 -4676 1352 -4642
rect 1266 -4710 1352 -4676
rect 1266 -4744 1292 -4710
rect 1326 -4744 1352 -4710
rect 1266 -4778 1352 -4744
rect 1266 -4812 1292 -4778
rect 1326 -4812 1352 -4778
rect 1266 -4846 1352 -4812
rect 1266 -4880 1292 -4846
rect 1326 -4880 1352 -4846
rect 1266 -4914 1352 -4880
rect 1266 -4948 1292 -4914
rect 1326 -4948 1352 -4914
rect 1266 -4982 1352 -4948
rect 1266 -5016 1292 -4982
rect 1326 -5016 1352 -4982
rect 1266 -5050 1352 -5016
rect 1266 -5084 1292 -5050
rect 1326 -5084 1352 -5050
rect 1266 -5118 1352 -5084
rect 1266 -5152 1292 -5118
rect 1326 -5152 1352 -5118
rect 1266 -5186 1352 -5152
rect 1266 -5220 1292 -5186
rect 1326 -5220 1352 -5186
rect 1266 -5254 1352 -5220
rect 1266 -5288 1292 -5254
rect 1326 -5288 1352 -5254
rect 1266 -5322 1352 -5288
rect 1266 -5356 1292 -5322
rect 1326 -5356 1352 -5322
rect 1266 -5384 1352 -5356
rect 2330 -4438 2416 -4384
rect 2330 -4472 2356 -4438
rect 2390 -4472 2416 -4438
rect 2330 -4506 2416 -4472
rect 2330 -4540 2356 -4506
rect 2390 -4540 2416 -4506
rect 2330 -4574 2416 -4540
rect 2330 -4608 2356 -4574
rect 2390 -4608 2416 -4574
rect 2330 -4642 2416 -4608
rect 2330 -4676 2356 -4642
rect 2390 -4676 2416 -4642
rect 2330 -4710 2416 -4676
rect 2330 -4744 2356 -4710
rect 2390 -4744 2416 -4710
rect 2330 -4778 2416 -4744
rect 2330 -4812 2356 -4778
rect 2390 -4812 2416 -4778
rect 2330 -4846 2416 -4812
rect 2330 -4880 2356 -4846
rect 2390 -4880 2416 -4846
rect 2330 -4914 2416 -4880
rect 2330 -4948 2356 -4914
rect 2390 -4948 2416 -4914
rect 2330 -4982 2416 -4948
rect 2330 -5016 2356 -4982
rect 2390 -5016 2416 -4982
rect 2330 -5050 2416 -5016
rect 2330 -5084 2356 -5050
rect 2390 -5084 2416 -5050
rect 2330 -5118 2416 -5084
rect 2330 -5152 2356 -5118
rect 2390 -5152 2416 -5118
rect 2330 -5186 2416 -5152
rect 2330 -5220 2356 -5186
rect 2390 -5220 2416 -5186
rect 2330 -5254 2416 -5220
rect 2330 -5288 2356 -5254
rect 2390 -5288 2416 -5254
rect 2330 -5322 2416 -5288
rect 2330 -5356 2356 -5322
rect 2390 -5356 2416 -5322
rect 2330 -5384 2416 -5356
<< nsubdiff >>
rect -4436 -1366 -4350 -1308
rect -4436 -1400 -4410 -1366
rect -4376 -1400 -4350 -1366
rect -4436 -1434 -4350 -1400
rect -4436 -1468 -4410 -1434
rect -4376 -1468 -4350 -1434
rect -4436 -1502 -4350 -1468
rect -4436 -1536 -4410 -1502
rect -4376 -1536 -4350 -1502
rect -4436 -1570 -4350 -1536
rect -4436 -1604 -4410 -1570
rect -4376 -1604 -4350 -1570
rect -4436 -1638 -4350 -1604
rect -4436 -1672 -4410 -1638
rect -4376 -1672 -4350 -1638
rect -4436 -1706 -4350 -1672
rect -4436 -1740 -4410 -1706
rect -4376 -1740 -4350 -1706
rect -4436 -1774 -4350 -1740
rect -4436 -1808 -4410 -1774
rect -4376 -1808 -4350 -1774
rect -4436 -1842 -4350 -1808
rect -4436 -1876 -4410 -1842
rect -4376 -1876 -4350 -1842
rect -4436 -1910 -4350 -1876
rect -4436 -1944 -4410 -1910
rect -4376 -1944 -4350 -1910
rect -4436 -1978 -4350 -1944
rect -4436 -2012 -4410 -1978
rect -4376 -2012 -4350 -1978
rect -4436 -2046 -4350 -2012
rect -4436 -2080 -4410 -2046
rect -4376 -2080 -4350 -2046
rect -4436 -2108 -4350 -2080
rect -304 -1362 -238 -1308
rect -304 -1396 -298 -1362
rect -264 -1396 -238 -1362
rect -304 -1430 -238 -1396
rect -304 -1464 -298 -1430
rect -264 -1464 -238 -1430
rect -304 -1498 -238 -1464
rect -304 -1532 -298 -1498
rect -264 -1532 -238 -1498
rect -304 -1566 -238 -1532
rect -304 -1600 -298 -1566
rect -264 -1600 -238 -1566
rect -304 -1634 -238 -1600
rect -304 -1668 -298 -1634
rect -264 -1668 -238 -1634
rect -304 -1702 -238 -1668
rect -304 -1736 -298 -1702
rect -264 -1736 -238 -1702
rect -304 -1770 -238 -1736
rect -304 -1804 -298 -1770
rect -264 -1804 -238 -1770
rect -304 -1838 -238 -1804
rect -304 -1872 -298 -1838
rect -264 -1872 -238 -1838
rect -304 -1906 -238 -1872
rect -304 -1940 -298 -1906
rect -264 -1940 -238 -1906
rect -304 -1974 -238 -1940
rect -304 -2008 -298 -1974
rect -264 -2008 -238 -1974
rect -304 -2042 -238 -2008
rect -304 -2076 -298 -2042
rect -264 -2076 -238 -2042
rect -304 -2110 -238 -2076
rect -304 -2144 -298 -2110
rect -264 -2144 -238 -2110
rect -304 -2178 -238 -2144
rect -304 -2212 -298 -2178
rect -264 -2212 -238 -2178
rect -304 -2246 -238 -2212
rect -304 -2280 -298 -2246
rect -264 -2280 -238 -2246
rect -304 -2308 -238 -2280
rect 740 -1362 826 -1308
rect 740 -1396 766 -1362
rect 800 -1396 826 -1362
rect 740 -1430 826 -1396
rect 740 -1464 766 -1430
rect 800 -1464 826 -1430
rect 740 -1498 826 -1464
rect 740 -1532 766 -1498
rect 800 -1532 826 -1498
rect 740 -1566 826 -1532
rect 740 -1600 766 -1566
rect 800 -1600 826 -1566
rect 740 -1634 826 -1600
rect 740 -1668 766 -1634
rect 800 -1668 826 -1634
rect 740 -1702 826 -1668
rect 740 -1736 766 -1702
rect 800 -1736 826 -1702
rect 740 -1770 826 -1736
rect 740 -1804 766 -1770
rect 800 -1804 826 -1770
rect 740 -1838 826 -1804
rect 740 -1872 766 -1838
rect 800 -1872 826 -1838
rect 740 -1906 826 -1872
rect 740 -1940 766 -1906
rect 800 -1940 826 -1906
rect 740 -1974 826 -1940
rect 740 -2008 766 -1974
rect 800 -2008 826 -1974
rect 740 -2042 826 -2008
rect 740 -2076 766 -2042
rect 800 -2076 826 -2042
rect 740 -2110 826 -2076
rect 740 -2144 766 -2110
rect 800 -2144 826 -2110
rect 740 -2178 826 -2144
rect 740 -2212 766 -2178
rect 800 -2212 826 -2178
rect 740 -2246 826 -2212
rect 740 -2280 766 -2246
rect 800 -2280 826 -2246
rect 740 -2308 826 -2280
rect 1804 -1362 1890 -1308
rect 1804 -1396 1830 -1362
rect 1864 -1396 1890 -1362
rect 1804 -1430 1890 -1396
rect 1804 -1464 1830 -1430
rect 1864 -1464 1890 -1430
rect 1804 -1498 1890 -1464
rect 1804 -1532 1830 -1498
rect 1864 -1532 1890 -1498
rect 1804 -1566 1890 -1532
rect 1804 -1600 1830 -1566
rect 1864 -1600 1890 -1566
rect 1804 -1634 1890 -1600
rect 1804 -1668 1830 -1634
rect 1864 -1668 1890 -1634
rect 1804 -1702 1890 -1668
rect 1804 -1736 1830 -1702
rect 1864 -1736 1890 -1702
rect 1804 -1770 1890 -1736
rect 1804 -1804 1830 -1770
rect 1864 -1804 1890 -1770
rect 1804 -1838 1890 -1804
rect 1804 -1872 1830 -1838
rect 1864 -1872 1890 -1838
rect 1804 -1906 1890 -1872
rect 1804 -1940 1830 -1906
rect 1864 -1940 1890 -1906
rect 1804 -1974 1890 -1940
rect 1804 -2008 1830 -1974
rect 1864 -2008 1890 -1974
rect 1804 -2042 1890 -2008
rect 1804 -2076 1830 -2042
rect 1864 -2076 1890 -2042
rect 1804 -2110 1890 -2076
rect 1804 -2144 1830 -2110
rect 1864 -2144 1890 -2110
rect 1804 -2178 1890 -2144
rect 1804 -2212 1830 -2178
rect 1864 -2212 1890 -2178
rect 1804 -2246 1890 -2212
rect 1804 -2280 1830 -2246
rect 1864 -2280 1890 -2246
rect 1804 -2308 1890 -2280
rect 2868 -1362 2954 -1308
rect 2868 -1396 2894 -1362
rect 2928 -1396 2954 -1362
rect 2868 -1430 2954 -1396
rect 2868 -1464 2894 -1430
rect 2928 -1464 2954 -1430
rect 2868 -1498 2954 -1464
rect 2868 -1532 2894 -1498
rect 2928 -1532 2954 -1498
rect 2868 -1566 2954 -1532
rect 2868 -1600 2894 -1566
rect 2928 -1600 2954 -1566
rect 2868 -1634 2954 -1600
rect 2868 -1668 2894 -1634
rect 2928 -1668 2954 -1634
rect 2868 -1702 2954 -1668
rect 2868 -1736 2894 -1702
rect 2928 -1736 2954 -1702
rect 2868 -1770 2954 -1736
rect 2868 -1804 2894 -1770
rect 2928 -1804 2954 -1770
rect 2868 -1838 2954 -1804
rect 2868 -1872 2894 -1838
rect 2928 -1872 2954 -1838
rect 2868 -1906 2954 -1872
rect 2868 -1940 2894 -1906
rect 2928 -1940 2954 -1906
rect 2868 -1974 2954 -1940
rect 2868 -2008 2894 -1974
rect 2928 -2008 2954 -1974
rect 2868 -2042 2954 -2008
rect 2868 -2076 2894 -2042
rect 2928 -2076 2954 -2042
rect 2868 -2110 2954 -2076
rect 2868 -2144 2894 -2110
rect 2928 -2144 2954 -2110
rect 2868 -2178 2954 -2144
rect 2868 -2212 2894 -2178
rect 2928 -2212 2954 -2178
rect 2868 -2246 2954 -2212
rect 2868 -2280 2894 -2246
rect 2928 -2280 2954 -2246
rect 2868 -2308 2954 -2280
rect 3932 -1362 3998 -1308
rect 3932 -1396 3958 -1362
rect 3992 -1396 3998 -1362
rect 3932 -1430 3998 -1396
rect 3932 -1464 3958 -1430
rect 3992 -1464 3998 -1430
rect 3932 -1498 3998 -1464
rect 3932 -1532 3958 -1498
rect 3992 -1532 3998 -1498
rect 3932 -1566 3998 -1532
rect 3932 -1600 3958 -1566
rect 3992 -1600 3998 -1566
rect 3932 -1634 3998 -1600
rect 3932 -1668 3958 -1634
rect 3992 -1668 3998 -1634
rect 3932 -1702 3998 -1668
rect 3932 -1736 3958 -1702
rect 3992 -1736 3998 -1702
rect 3932 -1770 3998 -1736
rect 3932 -1804 3958 -1770
rect 3992 -1804 3998 -1770
rect 3932 -1838 3998 -1804
rect 3932 -1872 3958 -1838
rect 3992 -1872 3998 -1838
rect 3932 -1906 3998 -1872
rect 3932 -1940 3958 -1906
rect 3992 -1940 3998 -1906
rect 3932 -1974 3998 -1940
rect 3932 -2008 3958 -1974
rect 3992 -2008 3998 -1974
rect 3932 -2042 3998 -2008
rect 3932 -2076 3958 -2042
rect 3992 -2076 3998 -2042
rect 3932 -2110 3998 -2076
rect 3932 -2144 3958 -2110
rect 3992 -2144 3998 -2110
rect 3932 -2178 3998 -2144
rect 3932 -2212 3958 -2178
rect 3992 -2212 3998 -2178
rect 3932 -2246 3998 -2212
rect 3932 -2280 3958 -2246
rect 3992 -2280 3998 -2246
rect 3932 -2308 3998 -2280
rect -2766 -4532 -2762 -4316
rect -2766 -4600 -2760 -4532
rect -2480 -4600 -2472 -4316
rect -1630 -4332 -1622 -4296
rect -1572 -4600 -1566 -4592
rect -1290 -4600 -1284 -4592
rect -2766 -4606 -2474 -4600
rect -1572 -4606 -1284 -4600
<< psubdiffcont >>
rect -3130 -1400 -3096 -1366
rect -3130 -1468 -3096 -1434
rect -3130 -1536 -3096 -1502
rect -3130 -1604 -3096 -1570
rect -3130 -1672 -3096 -1638
rect -3130 -1740 -3096 -1706
rect -3130 -1808 -3096 -1774
rect -3130 -1876 -3096 -1842
rect -3130 -1944 -3096 -1910
rect -3130 -2012 -3096 -1978
rect -3130 -2080 -3096 -2046
rect -2066 -1400 -2032 -1366
rect -2066 -1468 -2032 -1434
rect -2066 -1536 -2032 -1502
rect -2066 -1604 -2032 -1570
rect -2066 -1672 -2032 -1638
rect -2066 -1740 -2032 -1706
rect -2066 -1808 -2032 -1774
rect -2066 -1876 -2032 -1842
rect -2066 -1944 -2032 -1910
rect -2066 -2012 -2032 -1978
rect -2066 -2080 -2032 -2046
rect -1002 -1400 -968 -1366
rect -1002 -1468 -968 -1434
rect -1002 -1536 -968 -1502
rect -1002 -1604 -968 -1570
rect -1002 -1672 -968 -1638
rect -1002 -1740 -968 -1706
rect -1002 -1808 -968 -1774
rect -1002 -1876 -968 -1842
rect -1002 -1944 -968 -1910
rect -1002 -2012 -968 -1978
rect -1002 -2080 -968 -2046
rect -4410 -2954 -4376 -2920
rect -4410 -3022 -4376 -2988
rect -4410 -3090 -4376 -3056
rect -4410 -3158 -4376 -3124
rect -4410 -3226 -4376 -3192
rect -4410 -3294 -4376 -3260
rect -4410 -3362 -4376 -3328
rect -4410 -3430 -4376 -3396
rect -4410 -3498 -4376 -3464
rect -4410 -3566 -4376 -3532
rect -4410 -3634 -4376 -3600
rect -3130 -2954 -3096 -2920
rect -3130 -3022 -3096 -2988
rect -3130 -3090 -3096 -3056
rect -3130 -3158 -3096 -3124
rect -3130 -3226 -3096 -3192
rect -3130 -3294 -3096 -3260
rect -3130 -3362 -3096 -3328
rect -3130 -3430 -3096 -3396
rect -3130 -3498 -3096 -3464
rect -3130 -3566 -3096 -3532
rect -3130 -3634 -3096 -3600
rect -2066 -2954 -2032 -2920
rect -2066 -3022 -2032 -2988
rect -2066 -3090 -2032 -3056
rect -2066 -3158 -2032 -3124
rect -2066 -3226 -2032 -3192
rect -2066 -3294 -2032 -3260
rect -2066 -3362 -2032 -3328
rect -2066 -3430 -2032 -3396
rect -2066 -3498 -2032 -3464
rect -2066 -3566 -2032 -3532
rect -2066 -3634 -2032 -3600
rect -1002 -2954 -968 -2920
rect -1002 -3022 -968 -2988
rect -1002 -3090 -968 -3056
rect -1002 -3158 -968 -3124
rect -1002 -3226 -968 -3192
rect -1002 -3294 -968 -3260
rect -1002 -3362 -968 -3328
rect -1002 -3430 -968 -3396
rect -1002 -3498 -968 -3464
rect -1002 -3566 -968 -3532
rect -1002 -3634 -968 -3600
rect 2 -3024 36 -2990
rect 2 -3092 36 -3058
rect 2 -3160 36 -3126
rect 2 -3228 36 -3194
rect 2 -3296 36 -3262
rect 2 -3364 36 -3330
rect 2 -3432 36 -3398
rect 2 -3500 36 -3466
rect 2 -3568 36 -3534
rect 2 -3636 36 -3602
rect 2 -3704 36 -3670
rect 2 -3772 36 -3738
rect 2 -3840 36 -3806
rect 2 -3908 36 -3874
rect 466 -3024 500 -2990
rect 466 -3092 500 -3058
rect 466 -3160 500 -3126
rect 466 -3228 500 -3194
rect 466 -3296 500 -3262
rect 466 -3364 500 -3330
rect 466 -3432 500 -3398
rect 466 -3500 500 -3466
rect 466 -3568 500 -3534
rect 466 -3636 500 -3602
rect 466 -3704 500 -3670
rect 466 -3772 500 -3738
rect 466 -3840 500 -3806
rect 466 -3908 500 -3874
rect 1530 -3024 1564 -2990
rect 1530 -3092 1564 -3058
rect 1530 -3160 1564 -3126
rect 1530 -3228 1564 -3194
rect 1530 -3296 1564 -3262
rect 1530 -3364 1564 -3330
rect 1530 -3432 1564 -3398
rect 1530 -3500 1564 -3466
rect 1530 -3568 1564 -3534
rect 1530 -3636 1564 -3602
rect 1530 -3704 1564 -3670
rect 1530 -3772 1564 -3738
rect 1530 -3840 1564 -3806
rect 1530 -3908 1564 -3874
rect 2130 -3024 2164 -2990
rect 2130 -3092 2164 -3058
rect 2130 -3160 2164 -3126
rect 2130 -3228 2164 -3194
rect 2130 -3296 2164 -3262
rect 2130 -3364 2164 -3330
rect 2130 -3432 2164 -3398
rect 2130 -3500 2164 -3466
rect 2130 -3568 2164 -3534
rect 2130 -3636 2164 -3602
rect 2130 -3704 2164 -3670
rect 2130 -3772 2164 -3738
rect 2130 -3840 2164 -3806
rect 2130 -3908 2164 -3874
rect 2594 -3024 2628 -2990
rect 2594 -3092 2628 -3058
rect 2594 -3160 2628 -3126
rect 2594 -3228 2628 -3194
rect 2594 -3296 2628 -3262
rect 2594 -3364 2628 -3330
rect 2594 -3432 2628 -3398
rect 2594 -3500 2628 -3466
rect 2594 -3568 2628 -3534
rect 2594 -3636 2628 -3602
rect 2594 -3704 2628 -3670
rect 2594 -3772 2628 -3738
rect 2594 -3840 2628 -3806
rect 2594 -3908 2628 -3874
rect 3658 -3024 3692 -2990
rect 3658 -3092 3692 -3058
rect 3658 -3160 3692 -3126
rect 3658 -3228 3692 -3194
rect 3658 -3296 3692 -3262
rect 3658 -3364 3692 -3330
rect 3658 -3432 3692 -3398
rect 3658 -3500 3692 -3466
rect 3658 -3568 3692 -3534
rect 3658 -3636 3692 -3602
rect 3658 -3704 3692 -3670
rect 3658 -3772 3692 -3738
rect 3658 -3840 3692 -3806
rect 3658 -3908 3692 -3874
rect 1292 -4472 1326 -4438
rect 1292 -4540 1326 -4506
rect 1292 -4608 1326 -4574
rect 1292 -4676 1326 -4642
rect 1292 -4744 1326 -4710
rect 1292 -4812 1326 -4778
rect 1292 -4880 1326 -4846
rect 1292 -4948 1326 -4914
rect 1292 -5016 1326 -4982
rect 1292 -5084 1326 -5050
rect 1292 -5152 1326 -5118
rect 1292 -5220 1326 -5186
rect 1292 -5288 1326 -5254
rect 1292 -5356 1326 -5322
rect 2356 -4472 2390 -4438
rect 2356 -4540 2390 -4506
rect 2356 -4608 2390 -4574
rect 2356 -4676 2390 -4642
rect 2356 -4744 2390 -4710
rect 2356 -4812 2390 -4778
rect 2356 -4880 2390 -4846
rect 2356 -4948 2390 -4914
rect 2356 -5016 2390 -4982
rect 2356 -5084 2390 -5050
rect 2356 -5152 2390 -5118
rect 2356 -5220 2390 -5186
rect 2356 -5288 2390 -5254
rect 2356 -5356 2390 -5322
<< nsubdiffcont >>
rect -4410 -1400 -4376 -1366
rect -4410 -1468 -4376 -1434
rect -4410 -1536 -4376 -1502
rect -4410 -1604 -4376 -1570
rect -4410 -1672 -4376 -1638
rect -4410 -1740 -4376 -1706
rect -4410 -1808 -4376 -1774
rect -4410 -1876 -4376 -1842
rect -4410 -1944 -4376 -1910
rect -4410 -2012 -4376 -1978
rect -4410 -2080 -4376 -2046
rect -298 -1396 -264 -1362
rect -298 -1464 -264 -1430
rect -298 -1532 -264 -1498
rect -298 -1600 -264 -1566
rect -298 -1668 -264 -1634
rect -298 -1736 -264 -1702
rect -298 -1804 -264 -1770
rect -298 -1872 -264 -1838
rect -298 -1940 -264 -1906
rect -298 -2008 -264 -1974
rect -298 -2076 -264 -2042
rect -298 -2144 -264 -2110
rect -298 -2212 -264 -2178
rect -298 -2280 -264 -2246
rect 766 -1396 800 -1362
rect 766 -1464 800 -1430
rect 766 -1532 800 -1498
rect 766 -1600 800 -1566
rect 766 -1668 800 -1634
rect 766 -1736 800 -1702
rect 766 -1804 800 -1770
rect 766 -1872 800 -1838
rect 766 -1940 800 -1906
rect 766 -2008 800 -1974
rect 766 -2076 800 -2042
rect 766 -2144 800 -2110
rect 766 -2212 800 -2178
rect 766 -2280 800 -2246
rect 1830 -1396 1864 -1362
rect 1830 -1464 1864 -1430
rect 1830 -1532 1864 -1498
rect 1830 -1600 1864 -1566
rect 1830 -1668 1864 -1634
rect 1830 -1736 1864 -1702
rect 1830 -1804 1864 -1770
rect 1830 -1872 1864 -1838
rect 1830 -1940 1864 -1906
rect 1830 -2008 1864 -1974
rect 1830 -2076 1864 -2042
rect 1830 -2144 1864 -2110
rect 1830 -2212 1864 -2178
rect 1830 -2280 1864 -2246
rect 2894 -1396 2928 -1362
rect 2894 -1464 2928 -1430
rect 2894 -1532 2928 -1498
rect 2894 -1600 2928 -1566
rect 2894 -1668 2928 -1634
rect 2894 -1736 2928 -1702
rect 2894 -1804 2928 -1770
rect 2894 -1872 2928 -1838
rect 2894 -1940 2928 -1906
rect 2894 -2008 2928 -1974
rect 2894 -2076 2928 -2042
rect 2894 -2144 2928 -2110
rect 2894 -2212 2928 -2178
rect 2894 -2280 2928 -2246
rect 3958 -1396 3992 -1362
rect 3958 -1464 3992 -1430
rect 3958 -1532 3992 -1498
rect 3958 -1600 3992 -1566
rect 3958 -1668 3992 -1634
rect 3958 -1736 3992 -1702
rect 3958 -1804 3992 -1770
rect 3958 -1872 3992 -1838
rect 3958 -1940 3992 -1906
rect 3958 -2008 3992 -1974
rect 3958 -2076 3992 -2042
rect 3958 -2144 3992 -2110
rect 3958 -2212 3992 -2178
rect 3958 -2280 3992 -2246
<< poly >>
rect -3906 -2198 -3890 -2146
rect -4948 -2832 -4828 -2780
<< locali >>
rect -4410 -1320 -4376 -1304
rect -4410 -2112 -4376 -2096
rect -3130 -1320 -3096 -1304
rect -3130 -2112 -3096 -2096
rect -2066 -1320 -2032 -1304
rect -2066 -2112 -2032 -2096
rect -1002 -1320 -968 -1304
rect -1002 -2112 -968 -2096
rect -298 -1320 -264 -1304
rect -298 -2312 -264 -2296
rect 766 -1320 800 -1304
rect 766 -2312 800 -2296
rect 1830 -1320 1864 -1304
rect 1830 -2312 1864 -2296
rect 2894 -1320 2928 -1304
rect 2894 -2312 2928 -2296
rect 3958 -1320 3992 -1304
rect 3958 -2312 3992 -2296
rect -4410 -2874 -4376 -2858
rect -4410 -3666 -4376 -3650
rect -3130 -2874 -3096 -2858
rect -3130 -3666 -3096 -3650
rect -2066 -2874 -2032 -2858
rect -2066 -3666 -2032 -3650
rect -1002 -2874 -968 -2858
rect -1002 -3666 -968 -3650
rect 2 -2948 36 -2932
rect 2 -3940 36 -3924
rect 466 -2948 500 -2932
rect 466 -3940 500 -3924
rect 1530 -2948 1564 -2932
rect 1530 -3940 1564 -3924
rect 2130 -2948 2164 -2932
rect 2130 -3940 2164 -3924
rect 2594 -2948 2628 -2932
rect 2594 -3940 2628 -3924
rect 3658 -2948 3692 -2932
rect 3658 -3940 3692 -3924
rect -2766 -4532 -2762 -4316
rect -2766 -4600 -2760 -4532
rect -2480 -4600 -2474 -4316
rect -2766 -4606 -2474 -4600
rect -1572 -4600 -1566 -4592
rect -1290 -4600 -1284 -4592
rect -1572 -4606 -1284 -4600
rect 1292 -4396 1326 -4380
rect 1292 -5388 1326 -5372
rect 2356 -4396 2390 -4380
rect 2356 -5388 2390 -5372
<< viali >>
rect -4410 -1366 -4376 -1320
rect -4410 -1400 -4376 -1366
rect -4410 -1434 -4376 -1400
rect -4410 -1468 -4376 -1434
rect -4410 -1502 -4376 -1468
rect -4410 -1536 -4376 -1502
rect -4410 -1570 -4376 -1536
rect -4410 -1604 -4376 -1570
rect -4410 -1638 -4376 -1604
rect -4410 -1672 -4376 -1638
rect -4410 -1706 -4376 -1672
rect -4410 -1740 -4376 -1706
rect -4410 -1774 -4376 -1740
rect -4410 -1808 -4376 -1774
rect -4410 -1842 -4376 -1808
rect -4410 -1876 -4376 -1842
rect -4410 -1910 -4376 -1876
rect -4410 -1944 -4376 -1910
rect -4410 -1978 -4376 -1944
rect -4410 -2012 -4376 -1978
rect -4410 -2046 -4376 -2012
rect -4410 -2080 -4376 -2046
rect -4410 -2096 -4376 -2080
rect -3130 -1366 -3096 -1320
rect -3130 -1400 -3096 -1366
rect -3130 -1434 -3096 -1400
rect -3130 -1468 -3096 -1434
rect -3130 -1502 -3096 -1468
rect -3130 -1536 -3096 -1502
rect -3130 -1570 -3096 -1536
rect -3130 -1604 -3096 -1570
rect -3130 -1638 -3096 -1604
rect -3130 -1672 -3096 -1638
rect -3130 -1706 -3096 -1672
rect -3130 -1740 -3096 -1706
rect -3130 -1774 -3096 -1740
rect -3130 -1808 -3096 -1774
rect -3130 -1842 -3096 -1808
rect -3130 -1876 -3096 -1842
rect -3130 -1910 -3096 -1876
rect -3130 -1944 -3096 -1910
rect -3130 -1978 -3096 -1944
rect -3130 -2012 -3096 -1978
rect -3130 -2046 -3096 -2012
rect -3130 -2080 -3096 -2046
rect -3130 -2096 -3096 -2080
rect -2066 -1366 -2032 -1320
rect -2066 -1400 -2032 -1366
rect -2066 -1434 -2032 -1400
rect -2066 -1468 -2032 -1434
rect -2066 -1502 -2032 -1468
rect -2066 -1536 -2032 -1502
rect -2066 -1570 -2032 -1536
rect -2066 -1604 -2032 -1570
rect -2066 -1638 -2032 -1604
rect -2066 -1672 -2032 -1638
rect -2066 -1706 -2032 -1672
rect -2066 -1740 -2032 -1706
rect -2066 -1774 -2032 -1740
rect -2066 -1808 -2032 -1774
rect -2066 -1842 -2032 -1808
rect -2066 -1876 -2032 -1842
rect -2066 -1910 -2032 -1876
rect -2066 -1944 -2032 -1910
rect -2066 -1978 -2032 -1944
rect -2066 -2012 -2032 -1978
rect -2066 -2046 -2032 -2012
rect -2066 -2080 -2032 -2046
rect -2066 -2096 -2032 -2080
rect -1002 -1366 -968 -1320
rect -1002 -1400 -968 -1366
rect -1002 -1434 -968 -1400
rect -1002 -1468 -968 -1434
rect -1002 -1502 -968 -1468
rect -1002 -1536 -968 -1502
rect -1002 -1570 -968 -1536
rect -1002 -1604 -968 -1570
rect -1002 -1638 -968 -1604
rect -1002 -1672 -968 -1638
rect -1002 -1706 -968 -1672
rect -1002 -1740 -968 -1706
rect -1002 -1774 -968 -1740
rect -1002 -1808 -968 -1774
rect -1002 -1842 -968 -1808
rect -1002 -1876 -968 -1842
rect -1002 -1910 -968 -1876
rect -1002 -1944 -968 -1910
rect -1002 -1978 -968 -1944
rect -1002 -2012 -968 -1978
rect -1002 -2046 -968 -2012
rect -1002 -2080 -968 -2046
rect -1002 -2096 -968 -2080
rect -298 -1362 -264 -1320
rect -298 -1396 -264 -1362
rect -298 -1430 -264 -1396
rect -298 -1464 -264 -1430
rect -298 -1498 -264 -1464
rect -298 -1532 -264 -1498
rect -298 -1566 -264 -1532
rect -298 -1600 -264 -1566
rect -298 -1634 -264 -1600
rect -298 -1668 -264 -1634
rect -298 -1702 -264 -1668
rect -298 -1736 -264 -1702
rect -298 -1770 -264 -1736
rect -298 -1804 -264 -1770
rect -298 -1838 -264 -1804
rect -298 -1872 -264 -1838
rect -298 -1906 -264 -1872
rect -298 -1940 -264 -1906
rect -298 -1974 -264 -1940
rect -298 -2008 -264 -1974
rect -298 -2042 -264 -2008
rect -298 -2076 -264 -2042
rect -298 -2110 -264 -2076
rect -298 -2144 -264 -2110
rect -298 -2178 -264 -2144
rect -298 -2212 -264 -2178
rect -298 -2246 -264 -2212
rect -298 -2280 -264 -2246
rect -298 -2296 -264 -2280
rect 766 -1362 800 -1320
rect 766 -1396 800 -1362
rect 766 -1430 800 -1396
rect 766 -1464 800 -1430
rect 766 -1498 800 -1464
rect 766 -1532 800 -1498
rect 766 -1566 800 -1532
rect 766 -1600 800 -1566
rect 766 -1634 800 -1600
rect 766 -1668 800 -1634
rect 766 -1702 800 -1668
rect 766 -1736 800 -1702
rect 766 -1770 800 -1736
rect 766 -1804 800 -1770
rect 766 -1838 800 -1804
rect 766 -1872 800 -1838
rect 766 -1906 800 -1872
rect 766 -1940 800 -1906
rect 766 -1974 800 -1940
rect 766 -2008 800 -1974
rect 766 -2042 800 -2008
rect 766 -2076 800 -2042
rect 766 -2110 800 -2076
rect 766 -2144 800 -2110
rect 766 -2178 800 -2144
rect 766 -2212 800 -2178
rect 766 -2246 800 -2212
rect 766 -2280 800 -2246
rect 766 -2296 800 -2280
rect 1830 -1362 1864 -1320
rect 1830 -1396 1864 -1362
rect 1830 -1430 1864 -1396
rect 1830 -1464 1864 -1430
rect 1830 -1498 1864 -1464
rect 1830 -1532 1864 -1498
rect 1830 -1566 1864 -1532
rect 1830 -1600 1864 -1566
rect 1830 -1634 1864 -1600
rect 1830 -1668 1864 -1634
rect 1830 -1702 1864 -1668
rect 1830 -1736 1864 -1702
rect 1830 -1770 1864 -1736
rect 1830 -1804 1864 -1770
rect 1830 -1838 1864 -1804
rect 1830 -1872 1864 -1838
rect 1830 -1906 1864 -1872
rect 1830 -1940 1864 -1906
rect 1830 -1974 1864 -1940
rect 1830 -2008 1864 -1974
rect 1830 -2042 1864 -2008
rect 1830 -2076 1864 -2042
rect 1830 -2110 1864 -2076
rect 1830 -2144 1864 -2110
rect 1830 -2178 1864 -2144
rect 1830 -2212 1864 -2178
rect 1830 -2246 1864 -2212
rect 1830 -2280 1864 -2246
rect 1830 -2296 1864 -2280
rect 2894 -1362 2928 -1320
rect 2894 -1396 2928 -1362
rect 2894 -1430 2928 -1396
rect 2894 -1464 2928 -1430
rect 2894 -1498 2928 -1464
rect 2894 -1532 2928 -1498
rect 2894 -1566 2928 -1532
rect 2894 -1600 2928 -1566
rect 2894 -1634 2928 -1600
rect 2894 -1668 2928 -1634
rect 2894 -1702 2928 -1668
rect 2894 -1736 2928 -1702
rect 2894 -1770 2928 -1736
rect 2894 -1804 2928 -1770
rect 2894 -1838 2928 -1804
rect 2894 -1872 2928 -1838
rect 2894 -1906 2928 -1872
rect 2894 -1940 2928 -1906
rect 2894 -1974 2928 -1940
rect 2894 -2008 2928 -1974
rect 2894 -2042 2928 -2008
rect 2894 -2076 2928 -2042
rect 2894 -2110 2928 -2076
rect 2894 -2144 2928 -2110
rect 2894 -2178 2928 -2144
rect 2894 -2212 2928 -2178
rect 2894 -2246 2928 -2212
rect 2894 -2280 2928 -2246
rect 2894 -2296 2928 -2280
rect 3958 -1362 3992 -1320
rect 3958 -1396 3992 -1362
rect 3958 -1430 3992 -1396
rect 3958 -1464 3992 -1430
rect 3958 -1498 3992 -1464
rect 3958 -1532 3992 -1498
rect 3958 -1566 3992 -1532
rect 3958 -1600 3992 -1566
rect 3958 -1634 3992 -1600
rect 3958 -1668 3992 -1634
rect 3958 -1702 3992 -1668
rect 3958 -1736 3992 -1702
rect 3958 -1770 3992 -1736
rect 3958 -1804 3992 -1770
rect 3958 -1838 3992 -1804
rect 3958 -1872 3992 -1838
rect 3958 -1906 3992 -1872
rect 3958 -1940 3992 -1906
rect 3958 -1974 3992 -1940
rect 3958 -2008 3992 -1974
rect 3958 -2042 3992 -2008
rect 3958 -2076 3992 -2042
rect 3958 -2110 3992 -2076
rect 3958 -2144 3992 -2110
rect 3958 -2178 3992 -2144
rect 3958 -2212 3992 -2178
rect 3958 -2246 3992 -2212
rect 3958 -2280 3992 -2246
rect 3958 -2296 3992 -2280
rect -4410 -2920 -4376 -2874
rect -4410 -2954 -4376 -2920
rect -4410 -2988 -4376 -2954
rect -4410 -3022 -4376 -2988
rect -4410 -3056 -4376 -3022
rect -4410 -3090 -4376 -3056
rect -4410 -3124 -4376 -3090
rect -4410 -3158 -4376 -3124
rect -4410 -3192 -4376 -3158
rect -4410 -3226 -4376 -3192
rect -4410 -3260 -4376 -3226
rect -4410 -3294 -4376 -3260
rect -4410 -3328 -4376 -3294
rect -4410 -3362 -4376 -3328
rect -4410 -3396 -4376 -3362
rect -4410 -3430 -4376 -3396
rect -4410 -3464 -4376 -3430
rect -4410 -3498 -4376 -3464
rect -4410 -3532 -4376 -3498
rect -4410 -3566 -4376 -3532
rect -4410 -3600 -4376 -3566
rect -4410 -3634 -4376 -3600
rect -4410 -3650 -4376 -3634
rect -3130 -2920 -3096 -2874
rect -3130 -2954 -3096 -2920
rect -3130 -2988 -3096 -2954
rect -3130 -3022 -3096 -2988
rect -3130 -3056 -3096 -3022
rect -3130 -3090 -3096 -3056
rect -3130 -3124 -3096 -3090
rect -3130 -3158 -3096 -3124
rect -3130 -3192 -3096 -3158
rect -3130 -3226 -3096 -3192
rect -3130 -3260 -3096 -3226
rect -3130 -3294 -3096 -3260
rect -3130 -3328 -3096 -3294
rect -3130 -3362 -3096 -3328
rect -3130 -3396 -3096 -3362
rect -3130 -3430 -3096 -3396
rect -3130 -3464 -3096 -3430
rect -3130 -3498 -3096 -3464
rect -3130 -3532 -3096 -3498
rect -3130 -3566 -3096 -3532
rect -3130 -3600 -3096 -3566
rect -3130 -3634 -3096 -3600
rect -3130 -3650 -3096 -3634
rect -2066 -2920 -2032 -2874
rect -2066 -2954 -2032 -2920
rect -2066 -2988 -2032 -2954
rect -2066 -3022 -2032 -2988
rect -2066 -3056 -2032 -3022
rect -2066 -3090 -2032 -3056
rect -2066 -3124 -2032 -3090
rect -2066 -3158 -2032 -3124
rect -2066 -3192 -2032 -3158
rect -2066 -3226 -2032 -3192
rect -2066 -3260 -2032 -3226
rect -2066 -3294 -2032 -3260
rect -2066 -3328 -2032 -3294
rect -2066 -3362 -2032 -3328
rect -2066 -3396 -2032 -3362
rect -2066 -3430 -2032 -3396
rect -2066 -3464 -2032 -3430
rect -2066 -3498 -2032 -3464
rect -2066 -3532 -2032 -3498
rect -2066 -3566 -2032 -3532
rect -2066 -3600 -2032 -3566
rect -2066 -3634 -2032 -3600
rect -2066 -3650 -2032 -3634
rect -1002 -2920 -968 -2874
rect -1002 -2954 -968 -2920
rect -1002 -2988 -968 -2954
rect -1002 -3022 -968 -2988
rect -1002 -3056 -968 -3022
rect -1002 -3090 -968 -3056
rect -1002 -3124 -968 -3090
rect -1002 -3158 -968 -3124
rect -1002 -3192 -968 -3158
rect -1002 -3226 -968 -3192
rect -1002 -3260 -968 -3226
rect -1002 -3294 -968 -3260
rect -1002 -3328 -968 -3294
rect -1002 -3362 -968 -3328
rect -1002 -3396 -968 -3362
rect -1002 -3430 -968 -3396
rect -1002 -3464 -968 -3430
rect -1002 -3498 -968 -3464
rect -1002 -3532 -968 -3498
rect -1002 -3566 -968 -3532
rect -1002 -3600 -968 -3566
rect -1002 -3634 -968 -3600
rect -1002 -3650 -968 -3634
rect 2 -2990 36 -2948
rect 2 -3024 36 -2990
rect 2 -3058 36 -3024
rect 2 -3092 36 -3058
rect 2 -3126 36 -3092
rect 2 -3160 36 -3126
rect 2 -3194 36 -3160
rect 2 -3228 36 -3194
rect 2 -3262 36 -3228
rect 2 -3296 36 -3262
rect 2 -3330 36 -3296
rect 2 -3364 36 -3330
rect 2 -3398 36 -3364
rect 2 -3432 36 -3398
rect 2 -3466 36 -3432
rect 2 -3500 36 -3466
rect 2 -3534 36 -3500
rect 2 -3568 36 -3534
rect 2 -3602 36 -3568
rect 2 -3636 36 -3602
rect 2 -3670 36 -3636
rect 2 -3704 36 -3670
rect 2 -3738 36 -3704
rect 2 -3772 36 -3738
rect 2 -3806 36 -3772
rect 2 -3840 36 -3806
rect 2 -3874 36 -3840
rect 2 -3908 36 -3874
rect 2 -3924 36 -3908
rect 466 -2990 500 -2948
rect 466 -3024 500 -2990
rect 466 -3058 500 -3024
rect 466 -3092 500 -3058
rect 466 -3126 500 -3092
rect 466 -3160 500 -3126
rect 466 -3194 500 -3160
rect 466 -3228 500 -3194
rect 466 -3262 500 -3228
rect 466 -3296 500 -3262
rect 466 -3330 500 -3296
rect 466 -3364 500 -3330
rect 466 -3398 500 -3364
rect 466 -3432 500 -3398
rect 466 -3466 500 -3432
rect 466 -3500 500 -3466
rect 466 -3534 500 -3500
rect 466 -3568 500 -3534
rect 466 -3602 500 -3568
rect 466 -3636 500 -3602
rect 466 -3670 500 -3636
rect 466 -3704 500 -3670
rect 466 -3738 500 -3704
rect 466 -3772 500 -3738
rect 466 -3806 500 -3772
rect 466 -3840 500 -3806
rect 466 -3874 500 -3840
rect 466 -3908 500 -3874
rect 466 -3924 500 -3908
rect 1530 -2990 1564 -2948
rect 1530 -3024 1564 -2990
rect 1530 -3058 1564 -3024
rect 1530 -3092 1564 -3058
rect 1530 -3126 1564 -3092
rect 1530 -3160 1564 -3126
rect 1530 -3194 1564 -3160
rect 1530 -3228 1564 -3194
rect 1530 -3262 1564 -3228
rect 1530 -3296 1564 -3262
rect 1530 -3330 1564 -3296
rect 1530 -3364 1564 -3330
rect 1530 -3398 1564 -3364
rect 1530 -3432 1564 -3398
rect 1530 -3466 1564 -3432
rect 1530 -3500 1564 -3466
rect 1530 -3534 1564 -3500
rect 1530 -3568 1564 -3534
rect 1530 -3602 1564 -3568
rect 1530 -3636 1564 -3602
rect 1530 -3670 1564 -3636
rect 1530 -3704 1564 -3670
rect 1530 -3738 1564 -3704
rect 1530 -3772 1564 -3738
rect 1530 -3806 1564 -3772
rect 1530 -3840 1564 -3806
rect 1530 -3874 1564 -3840
rect 1530 -3908 1564 -3874
rect 1530 -3924 1564 -3908
rect 2130 -2990 2164 -2948
rect 2130 -3024 2164 -2990
rect 2130 -3058 2164 -3024
rect 2130 -3092 2164 -3058
rect 2130 -3126 2164 -3092
rect 2130 -3160 2164 -3126
rect 2130 -3194 2164 -3160
rect 2130 -3228 2164 -3194
rect 2130 -3262 2164 -3228
rect 2130 -3296 2164 -3262
rect 2130 -3330 2164 -3296
rect 2130 -3364 2164 -3330
rect 2130 -3398 2164 -3364
rect 2130 -3432 2164 -3398
rect 2130 -3466 2164 -3432
rect 2130 -3500 2164 -3466
rect 2130 -3534 2164 -3500
rect 2130 -3568 2164 -3534
rect 2130 -3602 2164 -3568
rect 2130 -3636 2164 -3602
rect 2130 -3670 2164 -3636
rect 2130 -3704 2164 -3670
rect 2130 -3738 2164 -3704
rect 2130 -3772 2164 -3738
rect 2130 -3806 2164 -3772
rect 2130 -3840 2164 -3806
rect 2130 -3874 2164 -3840
rect 2130 -3908 2164 -3874
rect 2130 -3924 2164 -3908
rect 2594 -2990 2628 -2948
rect 2594 -3024 2628 -2990
rect 2594 -3058 2628 -3024
rect 2594 -3092 2628 -3058
rect 2594 -3126 2628 -3092
rect 2594 -3160 2628 -3126
rect 2594 -3194 2628 -3160
rect 2594 -3228 2628 -3194
rect 2594 -3262 2628 -3228
rect 2594 -3296 2628 -3262
rect 2594 -3330 2628 -3296
rect 2594 -3364 2628 -3330
rect 2594 -3398 2628 -3364
rect 2594 -3432 2628 -3398
rect 2594 -3466 2628 -3432
rect 2594 -3500 2628 -3466
rect 2594 -3534 2628 -3500
rect 2594 -3568 2628 -3534
rect 2594 -3602 2628 -3568
rect 2594 -3636 2628 -3602
rect 2594 -3670 2628 -3636
rect 2594 -3704 2628 -3670
rect 2594 -3738 2628 -3704
rect 2594 -3772 2628 -3738
rect 2594 -3806 2628 -3772
rect 2594 -3840 2628 -3806
rect 2594 -3874 2628 -3840
rect 2594 -3908 2628 -3874
rect 2594 -3924 2628 -3908
rect 3658 -2990 3692 -2948
rect 3658 -3024 3692 -2990
rect 3658 -3058 3692 -3024
rect 3658 -3092 3692 -3058
rect 3658 -3126 3692 -3092
rect 3658 -3160 3692 -3126
rect 3658 -3194 3692 -3160
rect 3658 -3228 3692 -3194
rect 3658 -3262 3692 -3228
rect 3658 -3296 3692 -3262
rect 3658 -3330 3692 -3296
rect 3658 -3364 3692 -3330
rect 3658 -3398 3692 -3364
rect 3658 -3432 3692 -3398
rect 3658 -3466 3692 -3432
rect 3658 -3500 3692 -3466
rect 3658 -3534 3692 -3500
rect 3658 -3568 3692 -3534
rect 3658 -3602 3692 -3568
rect 3658 -3636 3692 -3602
rect 3658 -3670 3692 -3636
rect 3658 -3704 3692 -3670
rect 3658 -3738 3692 -3704
rect 3658 -3772 3692 -3738
rect 3658 -3806 3692 -3772
rect 3658 -3840 3692 -3806
rect 3658 -3874 3692 -3840
rect 3658 -3908 3692 -3874
rect 3658 -3924 3692 -3908
rect -2972 -4166 -2270 -4106
rect -2972 -4750 -2910 -4166
rect -2824 -4316 -2416 -4256
rect -2824 -4606 -2766 -4316
rect -2474 -4606 -2416 -4316
rect -2824 -4660 -2416 -4606
rect -2332 -4750 -2270 -4166
rect -2972 -4810 -2270 -4750
rect -1778 -4166 -1076 -4106
rect -1778 -4750 -1716 -4166
rect -1630 -4316 -1222 -4256
rect -1630 -4606 -1572 -4316
rect -1284 -4606 -1222 -4316
rect -1630 -4660 -1222 -4606
rect -1138 -4750 -1076 -4166
rect -1778 -4810 -1076 -4750
rect 1292 -4438 1326 -4396
rect 1292 -4472 1326 -4438
rect 1292 -4506 1326 -4472
rect 1292 -4540 1326 -4506
rect 1292 -4574 1326 -4540
rect 1292 -4608 1326 -4574
rect 1292 -4642 1326 -4608
rect 1292 -4676 1326 -4642
rect 1292 -4710 1326 -4676
rect 1292 -4744 1326 -4710
rect 1292 -4778 1326 -4744
rect 1292 -4812 1326 -4778
rect 1292 -4846 1326 -4812
rect 1292 -4880 1326 -4846
rect 1292 -4914 1326 -4880
rect 1292 -4948 1326 -4914
rect 1292 -4982 1326 -4948
rect 1292 -5016 1326 -4982
rect 1292 -5050 1326 -5016
rect 1292 -5084 1326 -5050
rect 1292 -5118 1326 -5084
rect 1292 -5152 1326 -5118
rect 1292 -5186 1326 -5152
rect 1292 -5220 1326 -5186
rect 1292 -5254 1326 -5220
rect 1292 -5288 1326 -5254
rect 1292 -5322 1326 -5288
rect 1292 -5356 1326 -5322
rect 1292 -5372 1326 -5356
rect 2356 -4438 2390 -4396
rect 2356 -4472 2390 -4438
rect 2356 -4506 2390 -4472
rect 2356 -4540 2390 -4506
rect 2356 -4574 2390 -4540
rect 2356 -4608 2390 -4574
rect 2356 -4642 2390 -4608
rect 2356 -4676 2390 -4642
rect 2356 -4710 2390 -4676
rect 2356 -4744 2390 -4710
rect 2356 -4778 2390 -4744
rect 2356 -4812 2390 -4778
rect 2356 -4846 2390 -4812
rect 2356 -4880 2390 -4846
rect 2356 -4914 2390 -4880
rect 2356 -4948 2390 -4914
rect 2356 -4982 2390 -4948
rect 2356 -5016 2390 -4982
rect 2356 -5050 2390 -5016
rect 2356 -5084 2390 -5050
rect 2356 -5118 2390 -5084
rect 2356 -5152 2390 -5118
rect 2356 -5186 2390 -5152
rect 2356 -5220 2390 -5186
rect 2356 -5254 2390 -5220
rect 2356 -5288 2390 -5254
rect 2356 -5322 2390 -5288
rect 2356 -5356 2390 -5322
rect 2356 -5372 2390 -5356
<< metal1 >>
rect -4490 -776 -4294 -770
rect -4950 -1320 -4898 -1314
rect -4950 -2078 -4898 -2072
rect -4490 -1320 -4294 -1226
rect -304 -776 -184 -770
rect -4490 -2096 -4410 -1320
rect -4376 -2096 -4294 -1320
rect -4490 -2108 -4294 -2096
rect -3866 -2146 -3710 -1308
rect -3672 -1320 -3616 -1308
rect -3224 -1320 -3172 -1314
rect -3136 -1320 -3090 -1308
rect -3054 -1318 -3002 -1312
rect -3672 -2072 -3670 -1320
rect -3618 -2072 -3616 -1320
rect -3672 -2138 -3616 -2072
rect -3226 -2096 -3224 -1320
rect -3172 -2096 -3170 -1320
rect -3226 -2106 -3170 -2096
rect -3136 -2096 -3130 -1320
rect -3096 -2096 -3090 -1320
rect -4886 -2198 -4880 -2146
rect -4512 -2198 -4506 -2146
rect -4280 -2198 -4274 -2146
rect -3726 -2198 -3710 -2146
rect -3680 -2190 -3674 -2138
rect -3232 -2190 -3226 -2138
rect -5400 -2832 -5356 -2780
rect -4512 -2832 -4506 -2780
rect -4280 -2832 -4274 -2780
rect -3906 -2832 -3900 -2780
rect -5400 -4252 -4896 -2832
rect -5400 -4356 -5356 -4252
rect -4902 -4356 -4896 -4252
rect -4490 -2874 -4296 -2862
rect -4490 -3650 -4410 -2874
rect -4376 -3650 -4296 -2874
rect -4490 -5426 -4296 -3650
rect -3866 -3662 -3710 -2198
rect -3136 -2874 -3090 -2096
rect -3056 -2096 -3054 -1318
rect -3002 -2096 -3000 -1318
rect -3056 -2102 -3000 -2096
rect -2606 -1320 -2554 -1314
rect -2606 -2102 -2554 -2096
rect -2162 -1318 -2106 -1312
rect -2162 -2090 -2160 -1318
rect -2108 -2090 -2106 -1318
rect -2162 -2100 -2106 -2090
rect -2072 -1320 -2026 -1308
rect -2072 -2096 -2066 -1320
rect -2032 -2096 -2026 -1320
rect -3000 -2190 -2994 -2138
rect -2626 -2190 -2620 -2138
rect -2542 -2190 -2536 -2138
rect -2168 -2190 -2162 -2138
rect -3000 -2780 -2626 -2190
rect -2536 -2780 -2162 -2190
rect -3000 -2832 -2994 -2780
rect -2626 -2832 -2620 -2780
rect -2542 -2832 -2536 -2780
rect -2168 -2832 -2162 -2780
rect -3136 -3650 -3130 -2874
rect -3096 -3650 -3090 -2874
rect -4490 -5882 -4296 -5876
rect -3136 -5420 -3090 -3650
rect -3056 -2874 -3000 -2864
rect -3056 -3650 -3054 -2874
rect -3002 -3650 -3000 -2874
rect -3056 -3656 -3000 -3650
rect -2606 -2874 -2554 -2868
rect -2162 -2874 -2106 -2864
rect -2162 -3646 -2160 -2874
rect -2108 -3646 -2106 -2874
rect -2072 -2874 -2026 -2096
rect -1992 -1318 -1936 -1312
rect -1992 -2096 -1990 -1318
rect -1938 -2096 -1936 -1318
rect -1992 -2106 -1936 -2096
rect -1542 -1320 -1490 -1314
rect -1542 -2102 -1490 -2096
rect -1098 -1318 -1042 -1312
rect -1098 -2090 -1096 -1318
rect -1044 -2090 -1042 -1318
rect -1098 -2100 -1042 -2090
rect -1008 -1320 -962 -1308
rect -1008 -2096 -1002 -1320
rect -968 -2096 -962 -1320
rect -1936 -2190 -1930 -2138
rect -1562 -2190 -1556 -2138
rect -1478 -2190 -1472 -2138
rect -1104 -2190 -1098 -2138
rect -1936 -2780 -1562 -2190
rect -1472 -2780 -1098 -2190
rect -1936 -2832 -1930 -2780
rect -1562 -2832 -1556 -2780
rect -1478 -2832 -1472 -2780
rect -1104 -2832 -1098 -2780
rect -2606 -3656 -2554 -3650
rect -2160 -3652 -2108 -3646
rect -2072 -3650 -2066 -2874
rect -2032 -3650 -2026 -2874
rect -1992 -2874 -1936 -2864
rect -1992 -3646 -1990 -2874
rect -1938 -3646 -1936 -2874
rect -1542 -2874 -1490 -2868
rect -2984 -4106 -2258 -4100
rect -2984 -4810 -2972 -4106
rect -2910 -4256 -2332 -4166
rect -2910 -4660 -2824 -4256
rect -2766 -4322 -2474 -4316
rect -2766 -4600 -2760 -4322
rect -2692 -4392 -2548 -4386
rect -2692 -4524 -2686 -4392
rect -2554 -4524 -2548 -4392
rect -2692 -4530 -2548 -4524
rect -2480 -4600 -2474 -4322
rect -2766 -4606 -2474 -4600
rect -2416 -4660 -2332 -4256
rect -2910 -4750 -2332 -4660
rect -2270 -4810 -2258 -4106
rect -3136 -5426 -3084 -5420
rect -3136 -5882 -3084 -5876
rect -2984 -5426 -2258 -4810
rect -2984 -5882 -2258 -5876
rect -2072 -5420 -2026 -3650
rect -1990 -3652 -1938 -3646
rect -1098 -2874 -1042 -2864
rect -1098 -3650 -1096 -2874
rect -1044 -3650 -1042 -2874
rect -1008 -2874 -962 -2096
rect -928 -1318 -872 -1312
rect -928 -2096 -926 -1318
rect -874 -2096 -872 -1318
rect -928 -2106 -872 -2096
rect -478 -1320 -426 -1314
rect -478 -2102 -426 -2096
rect -304 -1320 -184 -1226
rect 722 -776 842 -770
rect -872 -2190 -866 -2138
rect -498 -2190 -492 -2138
rect -872 -2780 -498 -2190
rect -304 -2296 -298 -1320
rect -264 -2296 -184 -1320
rect -304 -2308 -184 -2296
rect 224 -1320 276 -1314
rect 224 -2302 276 -2296
rect 722 -1320 842 -1226
rect 1786 -776 1906 -770
rect 722 -2296 766 -1320
rect 800 -2296 842 -1320
rect 722 -2308 842 -2296
rect 1286 -2346 1344 -1308
rect 1786 -1320 1906 -1226
rect 2850 -776 2970 -770
rect 1786 -2296 1830 -1320
rect 1864 -2296 1906 -1320
rect 1786 -2308 1906 -2296
rect 2350 -1320 2406 -1310
rect 2350 -2296 2352 -1320
rect 2404 -2296 2406 -1320
rect 2350 -2306 2406 -2296
rect 2850 -1320 2970 -1226
rect 3878 -776 3998 -770
rect 2850 -2296 2894 -1320
rect 2928 -2296 2970 -1320
rect 2850 -2308 2970 -2296
rect 3414 -2346 3472 -1308
rect 3878 -1320 3998 -1226
rect 3878 -2296 3958 -1320
rect 3992 -2296 3998 -1320
rect 3878 -2308 3998 -2296
rect -184 -2398 -178 -2346
rect 3916 -2398 3922 -2346
rect 126 -2534 132 -2430
rect 364 -2534 370 -2430
rect 2254 -2534 2260 -2430
rect 2492 -2534 2498 -2430
rect -230 -2678 -224 -2574
rect -120 -2678 -114 -2574
rect -224 -2718 -120 -2678
rect -872 -2832 -866 -2780
rect -498 -2832 -492 -2780
rect -230 -2822 -224 -2718
rect -120 -2822 -114 -2718
rect 132 -2854 370 -2534
rect 590 -2822 596 -2718
rect 1428 -2822 1434 -2718
rect -1008 -3650 -1002 -2874
rect -968 -3650 -962 -2874
rect -928 -2874 -872 -2864
rect -928 -3648 -926 -2874
rect -874 -3648 -872 -2874
rect -478 -2874 -426 -2868
rect -1542 -3656 -1490 -3650
rect -1096 -3656 -1044 -3650
rect -1790 -4106 -1064 -4100
rect -1790 -4810 -1778 -4106
rect -1716 -4256 -1138 -4166
rect -1716 -4660 -1630 -4256
rect -1572 -4322 -1284 -4316
rect -1572 -4600 -1566 -4322
rect -1498 -4392 -1354 -4386
rect -1498 -4524 -1492 -4392
rect -1360 -4524 -1354 -4392
rect -1498 -4530 -1354 -4524
rect -1290 -4600 -1284 -4322
rect -1572 -4606 -1284 -4600
rect -1222 -4660 -1138 -4256
rect -1716 -4750 -1138 -4660
rect -1076 -4810 -1064 -4106
rect -2072 -5426 -2020 -5420
rect -2072 -5882 -2020 -5876
rect -1790 -5426 -1064 -4810
rect -1790 -5882 -1064 -5876
rect -1008 -5420 -962 -3650
rect -926 -3654 -874 -3648
rect 132 -2906 138 -2854
rect 206 -2864 296 -2854
rect 206 -2906 212 -2864
rect 290 -2906 296 -2864
rect 364 -2906 370 -2854
rect 596 -2854 1434 -2822
rect 596 -2906 602 -2854
rect 970 -2866 1060 -2854
rect 970 -2906 976 -2866
rect 1054 -2906 1060 -2866
rect 1428 -2906 1434 -2854
rect 2260 -2854 2498 -2534
rect 4168 -2678 4174 -2574
rect 4336 -2678 4348 -2574
rect 2718 -2822 2724 -2718
rect 3556 -2822 3562 -2718
rect 2730 -2854 3556 -2822
rect 2260 -2906 2266 -2854
rect 2334 -2860 2424 -2854
rect 2334 -2906 2340 -2860
rect 2418 -2906 2424 -2860
rect 2492 -2906 2498 -2854
rect 2724 -2906 2730 -2854
rect 3098 -2866 3188 -2854
rect 3098 -2906 3104 -2866
rect 3182 -2906 3188 -2866
rect 3556 -2906 3562 -2854
rect -478 -3656 -426 -3650
rect -4 -2948 42 -2936
rect -4 -3924 2 -2948
rect 36 -3924 42 -2948
rect -4 -4108 42 -3924
rect 70 -3962 126 -2936
rect 222 -2948 278 -2938
rect 276 -3924 278 -2948
rect 222 -3934 278 -3924
rect 376 -3962 432 -2936
rect 70 -4066 76 -3962
rect 128 -4066 134 -3962
rect 368 -4066 374 -3962
rect 426 -4066 432 -3962
rect 460 -2948 506 -2936
rect 460 -3924 466 -2948
rect 500 -3924 506 -2948
rect 460 -4108 506 -3924
rect 534 -3962 590 -2936
rect 986 -2948 1042 -2938
rect 986 -3924 988 -2948
rect 1040 -3924 1042 -2948
rect 986 -3934 1042 -3924
rect 1440 -3962 1496 -2936
rect 534 -4066 540 -3962
rect 592 -4066 598 -3962
rect 722 -4066 728 -3962
rect 780 -4066 786 -3962
rect 1432 -4066 1438 -3962
rect 1490 -4066 1496 -3962
rect 1524 -2948 1570 -2936
rect 1524 -3924 1530 -2948
rect 1564 -3924 1570 -2948
rect -4 -4212 2 -4108
rect 54 -4212 60 -4108
rect 452 -4212 458 -4108
rect 510 -4212 516 -4108
rect 726 -4384 782 -4066
rect 1524 -4108 1570 -3924
rect 2124 -2948 2170 -2936
rect 2124 -3924 2130 -2948
rect 2164 -3924 2170 -2948
rect 2124 -4108 2170 -3924
rect 2198 -3962 2254 -2936
rect 2350 -2948 2406 -2938
rect 2404 -3924 2406 -2948
rect 2350 -3934 2406 -3924
rect 2504 -3962 2560 -2936
rect 2198 -4066 2204 -3962
rect 2256 -4066 2262 -3962
rect 2496 -4066 2502 -3962
rect 2554 -4066 2560 -3962
rect 2588 -2948 2634 -2936
rect 2588 -3924 2594 -2948
rect 2628 -3924 2634 -2948
rect 2588 -4108 2634 -3924
rect 2662 -3962 2718 -2936
rect 3114 -2948 3170 -2938
rect 3114 -3924 3116 -2948
rect 3168 -3924 3170 -2948
rect 3114 -3934 3170 -3924
rect 3568 -3962 3624 -2936
rect 2662 -4066 2668 -3962
rect 2720 -4066 2726 -3962
rect 2896 -4066 2902 -3962
rect 2954 -4066 2960 -3962
rect 3560 -4066 3566 -3962
rect 3618 -4066 3624 -3962
rect 3652 -2948 3698 -2936
rect 3652 -3924 3658 -2948
rect 3692 -3924 3698 -2948
rect 1278 -4212 1284 -4108
rect 1336 -4212 1342 -4108
rect 1516 -4212 1522 -4108
rect 1574 -4212 1580 -4108
rect 2116 -4212 2122 -4108
rect 2174 -4212 2180 -4108
rect 2342 -4212 2348 -4108
rect 2400 -4212 2406 -4108
rect 2580 -4212 2586 -4108
rect 2638 -4212 2644 -4108
rect 816 -4356 822 -4304
rect 1190 -4356 1196 -4304
rect 1286 -4384 1332 -4212
rect 1422 -4356 1428 -4304
rect 1796 -4356 1802 -4304
rect 1880 -4356 1886 -4304
rect 2254 -4356 2260 -4304
rect 2350 -4384 2396 -4212
rect 2486 -4356 2492 -4304
rect 2860 -4356 2866 -4304
rect 2900 -4384 2956 -4066
rect 3652 -4108 3698 -3924
rect 3634 -4212 3640 -4108
rect 3692 -4212 3698 -4108
rect 726 -5384 800 -4384
rect 1212 -4396 1406 -4384
rect 1212 -5372 1292 -4396
rect 1326 -5372 1406 -4396
rect 1212 -5384 1406 -5372
rect 1812 -4394 1868 -4384
rect 1812 -5370 1814 -4394
rect 1866 -5370 1868 -4394
rect 1812 -5380 1868 -5370
rect 2276 -4396 2470 -4384
rect 2276 -5372 2356 -4396
rect 2390 -5372 2470 -4396
rect 2276 -5384 2470 -5372
rect 2882 -5384 2956 -4384
rect 4174 -4992 4348 -2678
rect -1008 -5426 -956 -5420
rect -1008 -5882 -956 -5876
rect 1248 -5426 1368 -5384
rect 1248 -5882 1368 -5876
rect 2312 -5426 2432 -5384
rect 2312 -5882 2432 -5876
<< via1 >>
rect -4490 -1226 -4294 -776
rect -4950 -2072 -4898 -1320
rect -304 -1226 -184 -776
rect -3670 -2072 -3618 -1320
rect -3224 -2096 -3172 -1320
rect -4880 -2198 -4512 -2146
rect -4274 -2198 -3726 -2146
rect -3674 -2190 -3232 -2138
rect -5356 -2832 -4512 -2780
rect -4274 -2832 -3906 -2780
rect -5356 -4356 -4902 -4252
rect -3054 -2096 -3002 -1318
rect -2606 -2096 -2554 -1320
rect -2160 -2090 -2108 -1318
rect -2994 -2190 -2626 -2138
rect -2536 -2190 -2168 -2138
rect -2994 -2832 -2626 -2780
rect -2536 -2832 -2168 -2780
rect -4490 -5876 -4296 -5426
rect -3054 -3650 -3002 -2874
rect -2606 -3650 -2554 -2874
rect -2160 -3646 -2108 -2874
rect -1990 -2096 -1938 -1318
rect -1542 -2096 -1490 -1320
rect -1096 -2090 -1044 -1318
rect -1930 -2190 -1562 -2138
rect -1472 -2190 -1104 -2138
rect -1930 -2832 -1562 -2780
rect -1472 -2832 -1104 -2780
rect -1990 -3646 -1938 -2874
rect -2686 -4524 -2554 -4392
rect -3136 -5876 -3084 -5426
rect -2984 -5876 -2258 -5426
rect -1542 -3650 -1490 -2874
rect -1096 -3650 -1044 -2874
rect -926 -2096 -874 -1318
rect -478 -2096 -426 -1320
rect 722 -1226 842 -776
rect -866 -2190 -498 -2138
rect 224 -2296 276 -1320
rect 1786 -1226 1906 -776
rect 2850 -1226 2970 -776
rect 2352 -2296 2404 -1320
rect 3878 -1226 3998 -776
rect -178 -2398 3916 -2346
rect 132 -2534 364 -2430
rect 2260 -2534 2492 -2430
rect -224 -2678 -120 -2574
rect -866 -2832 -498 -2780
rect -224 -2822 -120 -2718
rect 596 -2822 1428 -2718
rect -926 -3648 -874 -2874
rect -1492 -4524 -1360 -4392
rect -2072 -5876 -2020 -5426
rect -1790 -5876 -1064 -5426
rect -478 -3650 -426 -2874
rect 138 -2906 206 -2854
rect 296 -2906 364 -2854
rect 602 -2906 970 -2854
rect 1060 -2906 1428 -2854
rect 4174 -2678 4336 -2574
rect 2724 -2822 3556 -2718
rect 2266 -2906 2334 -2854
rect 2424 -2906 2492 -2854
rect 2730 -2906 3098 -2854
rect 3188 -2906 3556 -2854
rect 222 -3924 276 -2948
rect 76 -4066 128 -3962
rect 374 -4066 426 -3962
rect 988 -3924 1040 -2948
rect 540 -4066 592 -3962
rect 728 -4066 780 -3962
rect 1438 -4066 1490 -3962
rect 2 -4212 54 -4108
rect 458 -4212 510 -4108
rect 2350 -3924 2404 -2948
rect 2204 -4066 2256 -3962
rect 2502 -4066 2554 -3962
rect 3116 -3924 3168 -2948
rect 2668 -4066 2720 -3962
rect 2902 -4066 2954 -3962
rect 3566 -4066 3618 -3962
rect 1284 -4212 1336 -4108
rect 1522 -4212 1574 -4108
rect 2122 -4212 2174 -4108
rect 2348 -4212 2400 -4108
rect 2586 -4212 2638 -4108
rect 822 -4356 1190 -4304
rect 1428 -4356 1796 -4304
rect 1886 -4356 2254 -4304
rect 2492 -4356 2860 -4304
rect 3640 -4212 3692 -4108
rect 1814 -5370 1866 -4394
rect -1008 -5876 -956 -5426
rect 1248 -5876 1368 -5426
rect 2312 -5876 2432 -5426
<< metal2 >>
rect -5400 -776 4348 -764
rect -5400 -1226 -4490 -776
rect -4294 -780 -304 -776
rect -4294 -1222 -2608 -780
rect -2552 -1222 -1544 -780
rect -1488 -1222 -480 -780
rect -424 -1222 -304 -780
rect -4294 -1226 -304 -1222
rect -184 -1226 722 -776
rect 842 -1226 1786 -776
rect 1906 -1226 2850 -776
rect 2970 -1226 3878 -776
rect 3998 -1226 4348 -776
rect -5400 -1232 4348 -1226
rect -4950 -1320 -3618 -1314
rect -4898 -2072 -3670 -1320
rect -4950 -2078 -3618 -2072
rect -3226 -1320 -3170 -1310
rect -3226 -2106 -3170 -2096
rect -3056 -1318 -3000 -1308
rect -3056 -2106 -3000 -2096
rect -2608 -1320 -2552 -1310
rect -2608 -2106 -2552 -2096
rect -2162 -1318 -2106 -1308
rect -2162 -2100 -2106 -2090
rect -1992 -1318 -1936 -1308
rect -1992 -2106 -1936 -2096
rect -1544 -1320 -1488 -1310
rect -1544 -2106 -1488 -2096
rect -1098 -1318 -1042 -1308
rect -1098 -2100 -1042 -2090
rect -928 -1318 -872 -1308
rect -928 -2106 -872 -2096
rect -480 -1320 -424 -1310
rect -480 -2106 -424 -2096
rect 222 -1320 278 -1310
rect -3680 -2138 -486 -2134
rect -4886 -2198 -4880 -2146
rect -4512 -2198 -4274 -2146
rect -3726 -2198 -3720 -2146
rect -3680 -2190 -3674 -2138
rect -3232 -2190 -2994 -2138
rect -2626 -2190 -2536 -2138
rect -2168 -2190 -1930 -2138
rect -1562 -2190 -1472 -2138
rect -1104 -2190 -866 -2138
rect -498 -2190 -486 -2138
rect -3680 -2194 -486 -2190
rect 222 -2306 278 -2296
rect 2350 -1320 2406 -1310
rect 2350 -2306 2406 -2296
rect -184 -2344 3112 -2342
rect -184 -2346 984 -2344
rect 1044 -2346 3112 -2344
rect 3172 -2346 3922 -2342
rect -184 -2398 -178 -2346
rect 3916 -2398 3922 -2346
rect -184 -2400 984 -2398
rect 1044 -2400 3922 -2398
rect -184 -2402 3922 -2400
rect -3066 -2436 132 -2430
rect -3066 -2528 -3056 -2436
rect -3000 -2528 -2162 -2436
rect -2106 -2528 -1992 -2436
rect -1936 -2528 -1098 -2436
rect -1042 -2528 -928 -2436
rect -872 -2528 132 -2436
rect -3066 -2534 132 -2528
rect 364 -2534 2260 -2430
rect 2492 -2534 2498 -2430
rect -3236 -2580 -224 -2574
rect -3236 -2672 -3226 -2580
rect -3170 -2672 -224 -2580
rect -3236 -2678 -224 -2672
rect -120 -2678 -114 -2574
rect 212 -2580 4174 -2574
rect 212 -2672 222 -2580
rect 278 -2672 2350 -2580
rect 2406 -2672 4174 -2580
rect 212 -2678 4174 -2672
rect 4336 -2678 4342 -2574
rect -3006 -2780 -486 -2776
rect -5362 -2832 -5356 -2780
rect -4512 -2832 -4274 -2780
rect -3906 -2832 -3900 -2780
rect -3006 -2832 -2994 -2780
rect -2626 -2832 -2536 -2780
rect -2168 -2832 -1930 -2780
rect -1562 -2832 -1472 -2780
rect -1104 -2832 -866 -2780
rect -498 -2832 -486 -2780
rect -230 -2822 -224 -2718
rect -120 -2822 596 -2718
rect 1428 -2822 2724 -2718
rect 3556 -2822 3562 -2718
rect -3006 -2836 -486 -2832
rect 132 -2854 370 -2850
rect -3056 -2874 -3000 -2864
rect -3056 -3660 -3000 -3650
rect -2608 -2874 -2552 -2864
rect -2608 -3660 -2552 -3650
rect -2162 -2874 -2106 -2864
rect -2162 -3656 -2106 -3646
rect -1992 -2874 -1936 -2864
rect -1992 -3656 -1936 -3646
rect -1544 -2874 -1488 -2864
rect -1544 -3660 -1488 -3650
rect -1098 -2874 -1042 -2864
rect -1098 -3660 -1042 -3650
rect -928 -2874 -872 -2864
rect -928 -3658 -872 -3648
rect -480 -2874 -424 -2864
rect 132 -2906 138 -2854
rect 206 -2906 296 -2854
rect 364 -2906 370 -2854
rect 132 -2910 370 -2906
rect 596 -2854 1434 -2850
rect 596 -2906 602 -2854
rect 970 -2906 1060 -2854
rect 1428 -2906 1434 -2854
rect 596 -2910 1434 -2906
rect 2260 -2854 2498 -2850
rect 2260 -2906 2266 -2854
rect 2334 -2906 2424 -2854
rect 2492 -2906 2498 -2854
rect 2260 -2910 2498 -2906
rect 2724 -2854 3562 -2850
rect 2724 -2906 2730 -2854
rect 3098 -2906 3188 -2854
rect 3556 -2906 3562 -2854
rect 2724 -2910 3562 -2906
rect -480 -3660 -424 -3650
rect 222 -2948 278 -2938
rect 222 -3934 278 -3924
rect 986 -2948 1042 -2938
rect 986 -3934 1042 -3924
rect 2350 -2948 2406 -2938
rect 2350 -3934 2406 -3924
rect 3114 -2948 3170 -2938
rect 3114 -3934 3170 -3924
rect 70 -4066 76 -3962
rect 128 -4066 374 -3962
rect 426 -4066 540 -3962
rect 592 -4066 728 -3962
rect 780 -4066 1438 -3962
rect 1490 -3968 2204 -3962
rect 1490 -4060 1812 -3968
rect 1868 -4060 2204 -3968
rect 1490 -4066 2204 -4060
rect 2256 -4066 2502 -3962
rect 2554 -4066 2668 -3962
rect 2720 -4066 2902 -3962
rect 2954 -4066 3566 -3962
rect 3618 -4066 3624 -3962
rect -4 -4212 2 -4108
rect 54 -4212 458 -4108
rect 510 -4212 1284 -4108
rect 1336 -4212 1522 -4108
rect 1574 -4212 2122 -4108
rect 2174 -4212 2348 -4108
rect 2400 -4212 2586 -4108
rect 2638 -4212 3640 -4108
rect 3692 -4212 3698 -4108
rect -5362 -4356 -5356 -4252
rect -4902 -4304 2866 -4252
rect -4902 -4356 822 -4304
rect 1190 -4356 1428 -4304
rect 1796 -4356 1886 -4304
rect 2254 -4356 2492 -4304
rect 2860 -4356 2866 -4304
rect -2692 -4392 -2548 -4386
rect -1498 -4392 -1354 -4386
rect -3232 -4402 -2686 -4392
rect -3232 -4514 -3222 -4402
rect -3166 -4514 -2686 -4402
rect -3232 -4524 -2686 -4514
rect -2554 -4524 -2548 -4392
rect -1998 -4402 -1492 -4392
rect -1998 -4514 -1988 -4402
rect -1932 -4514 -1492 -4402
rect -1998 -4524 -1492 -4514
rect -1360 -4524 -1354 -4392
rect -2692 -4530 -2548 -4524
rect -1498 -4530 -1354 -4524
rect 1812 -4394 1868 -4384
rect 1812 -5380 1868 -5370
rect -5400 -5426 4348 -5420
rect -5400 -5876 -4490 -5426
rect -4296 -5876 -3136 -5426
rect -3084 -5876 -2984 -5426
rect -2258 -5876 -2072 -5426
rect -2020 -5876 -1790 -5426
rect -1064 -5876 -1008 -5426
rect -956 -5876 1248 -5426
rect 1368 -5876 2312 -5426
rect 2432 -5876 4348 -5426
rect -5400 -5888 4348 -5876
<< via2 >>
rect -2608 -1222 -2552 -780
rect -1544 -1222 -1488 -780
rect -480 -1222 -424 -780
rect -3226 -2096 -3224 -1320
rect -3224 -2096 -3172 -1320
rect -3172 -2096 -3170 -1320
rect -3056 -2096 -3054 -1318
rect -3054 -2096 -3002 -1318
rect -3002 -2096 -3000 -1318
rect -2608 -2096 -2606 -1320
rect -2606 -2096 -2554 -1320
rect -2554 -2096 -2552 -1320
rect -2162 -2090 -2160 -1318
rect -2160 -2090 -2108 -1318
rect -2108 -2090 -2106 -1318
rect -1992 -2096 -1990 -1318
rect -1990 -2096 -1938 -1318
rect -1938 -2096 -1936 -1318
rect -1544 -2096 -1542 -1320
rect -1542 -2096 -1490 -1320
rect -1490 -2096 -1488 -1320
rect -1098 -2090 -1096 -1318
rect -1096 -2090 -1044 -1318
rect -1044 -2090 -1042 -1318
rect -928 -2096 -926 -1318
rect -926 -2096 -874 -1318
rect -874 -2096 -872 -1318
rect -480 -2096 -478 -1320
rect -478 -2096 -426 -1320
rect -426 -2096 -424 -1320
rect 222 -2296 224 -1320
rect 224 -2296 276 -1320
rect 276 -2296 278 -1320
rect 2350 -2296 2352 -1320
rect 2352 -2296 2404 -1320
rect 2404 -2296 2406 -1320
rect 984 -2346 1044 -2344
rect 3112 -2346 3172 -2342
rect 984 -2398 1044 -2346
rect 3112 -2398 3172 -2346
rect 984 -2400 1044 -2398
rect -3056 -2528 -3000 -2436
rect -2162 -2528 -2106 -2436
rect -1992 -2528 -1936 -2436
rect -1098 -2528 -1042 -2436
rect -928 -2528 -872 -2436
rect -3226 -2672 -3170 -2580
rect 222 -2672 278 -2580
rect 2350 -2672 2406 -2580
rect -3056 -3650 -3054 -2874
rect -3054 -3650 -3002 -2874
rect -3002 -3650 -3000 -2874
rect -2608 -3650 -2606 -2874
rect -2606 -3650 -2554 -2874
rect -2554 -3650 -2552 -2874
rect -2162 -3646 -2160 -2874
rect -2160 -3646 -2108 -2874
rect -2108 -3646 -2106 -2874
rect -1992 -3646 -1990 -2874
rect -1990 -3646 -1938 -2874
rect -1938 -3646 -1936 -2874
rect -1544 -3650 -1542 -2874
rect -1542 -3650 -1490 -2874
rect -1490 -3650 -1488 -2874
rect -1098 -3650 -1096 -2874
rect -1096 -3650 -1044 -2874
rect -1044 -3650 -1042 -2874
rect -928 -3648 -926 -2874
rect -926 -3648 -874 -2874
rect -874 -3648 -872 -2874
rect -480 -3650 -478 -2874
rect -478 -3650 -426 -2874
rect -426 -3650 -424 -2874
rect 222 -3924 276 -2948
rect 276 -3924 278 -2948
rect 986 -3924 988 -2948
rect 988 -3924 1040 -2948
rect 1040 -3924 1042 -2948
rect 2350 -3924 2404 -2948
rect 2404 -3924 2406 -2948
rect 3114 -3924 3116 -2948
rect 3116 -3924 3168 -2948
rect 3168 -3924 3170 -2948
rect 1812 -4060 1868 -3968
rect -3222 -4514 -3166 -4402
rect -1988 -4514 -1932 -4402
rect 1812 -5370 1814 -4394
rect 1814 -5370 1866 -4394
rect 1866 -5370 1868 -4394
<< metal3 >>
rect -2614 -780 -2546 -770
rect -2614 -1222 -2608 -780
rect -2552 -1222 -2546 -780
rect -3232 -1320 -3164 -1314
rect -3232 -2096 -3226 -1320
rect -3170 -2096 -3164 -1320
rect -3232 -2580 -3164 -2096
rect -3232 -2672 -3226 -2580
rect -3170 -2672 -3164 -2580
rect -3232 -4392 -3164 -2672
rect -3062 -1318 -2994 -1312
rect -3062 -2096 -3056 -1318
rect -3000 -2096 -2994 -1318
rect -3062 -2436 -2994 -2096
rect -3062 -2528 -3056 -2436
rect -3000 -2528 -2994 -2436
rect -3062 -2874 -2994 -2528
rect -3062 -3650 -3056 -2874
rect -3000 -3650 -2994 -2874
rect -3062 -3656 -2994 -3650
rect -2614 -1320 -2546 -1222
rect -1550 -780 -1482 -770
rect -1550 -1222 -1544 -780
rect -1488 -1222 -1482 -780
rect -2614 -2096 -2608 -1320
rect -2552 -2096 -2546 -1320
rect -2614 -2874 -2546 -2096
rect -2614 -3650 -2608 -2874
rect -2552 -3650 -2546 -2874
rect -2614 -3656 -2546 -3650
rect -2168 -1318 -2100 -1312
rect -2168 -2090 -2162 -1318
rect -2106 -2090 -2100 -1318
rect -2168 -2436 -2100 -2090
rect -2168 -2528 -2162 -2436
rect -2106 -2528 -2100 -2436
rect -2168 -2874 -2100 -2528
rect -2168 -3646 -2162 -2874
rect -2106 -3646 -2100 -2874
rect -2168 -3652 -2100 -3646
rect -1998 -1318 -1930 -1312
rect -1998 -2096 -1992 -1318
rect -1936 -2096 -1930 -1318
rect -1998 -2436 -1930 -2096
rect -1998 -2528 -1992 -2436
rect -1936 -2528 -1930 -2436
rect -1998 -2874 -1930 -2528
rect -1998 -3646 -1992 -2874
rect -1936 -3646 -1930 -2874
rect -1998 -4392 -1930 -3646
rect -1550 -1320 -1482 -1222
rect -486 -780 -418 -770
rect -486 -1222 -480 -780
rect -424 -1222 -418 -780
rect -1550 -2096 -1544 -1320
rect -1488 -2096 -1482 -1320
rect -1550 -2874 -1482 -2096
rect -1550 -3650 -1544 -2874
rect -1488 -3650 -1482 -2874
rect -1550 -3656 -1482 -3650
rect -1104 -1318 -1036 -1312
rect -1104 -2090 -1098 -1318
rect -1042 -2090 -1036 -1318
rect -1104 -2436 -1036 -2090
rect -1104 -2528 -1098 -2436
rect -1042 -2528 -1036 -2436
rect -1104 -2874 -1036 -2528
rect -1104 -3650 -1098 -2874
rect -1042 -3650 -1036 -2874
rect -1104 -3656 -1036 -3650
rect -934 -1318 -866 -1312
rect -934 -2096 -928 -1318
rect -872 -2096 -866 -1318
rect -934 -2436 -866 -2096
rect -934 -2528 -928 -2436
rect -872 -2528 -866 -2436
rect -934 -2874 -866 -2528
rect -934 -3648 -928 -2874
rect -872 -3648 -866 -2874
rect -934 -3654 -866 -3648
rect -486 -1320 -418 -1222
rect -486 -2096 -480 -1320
rect -424 -2096 -418 -1320
rect -486 -2874 -418 -2096
rect -486 -3650 -480 -2874
rect -424 -3650 -418 -2874
rect -486 -3656 -418 -3650
rect 216 -1320 284 -1314
rect 216 -2296 222 -1320
rect 278 -2296 284 -1320
rect 216 -2580 284 -2296
rect 2344 -1320 2412 -1314
rect 2344 -2296 2350 -1320
rect 2406 -2296 2412 -1320
rect 978 -2344 1050 -2338
rect 978 -2400 984 -2344
rect 1044 -2400 1050 -2344
rect 978 -2406 1050 -2400
rect 216 -2672 222 -2580
rect 278 -2672 284 -2580
rect 216 -2948 284 -2672
rect 216 -3924 222 -2948
rect 278 -3924 284 -2948
rect 216 -3930 284 -3924
rect 980 -2948 1048 -2406
rect 980 -3924 986 -2948
rect 1042 -3924 1048 -2948
rect 980 -3930 1048 -3924
rect 2344 -2580 2412 -2296
rect 3106 -2342 3178 -2336
rect 3106 -2398 3112 -2342
rect 3172 -2398 3178 -2342
rect 3106 -2404 3178 -2398
rect 2344 -2672 2350 -2580
rect 2406 -2672 2412 -2580
rect 2344 -2948 2412 -2672
rect 2344 -3924 2350 -2948
rect 2406 -3924 2412 -2948
rect 2344 -3930 2412 -3924
rect 3108 -2948 3176 -2404
rect 3108 -3924 3114 -2948
rect 3170 -3924 3176 -2948
rect 3108 -3930 3176 -3924
rect 1806 -3968 1874 -3962
rect 1806 -4060 1812 -3968
rect 1868 -4060 1874 -3968
rect -3232 -4402 -3160 -4392
rect -3232 -4514 -3222 -4402
rect -3166 -4514 -3160 -4402
rect -3232 -4524 -3160 -4514
rect -1998 -4402 -1926 -4392
rect -1998 -4514 -1988 -4402
rect -1932 -4514 -1926 -4402
rect -1998 -4524 -1926 -4514
rect 1806 -4394 1874 -4060
rect 1806 -5370 1812 -4394
rect 1868 -5370 1874 -4394
rect 1806 -5376 1874 -5370
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M1
timestamp 1681340463
transform -1 0 -4696 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M2
timestamp 1681340463
transform 1 0 -4090 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__pfet_01v8_lvt_HLT7ZV  M3
timestamp 1681340463
transform 1 0 -4090 0 1 -1744
box -294 -464 294 498
use sky130_fd_pr__pfet_01v8_lvt_HLT7ZV  M4
timestamp 1681340463
transform -1 0 -4696 0 1 -1744
box -294 -464 294 498
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M5
timestamp 1681340463
transform -1 0 -3416 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M61
timestamp 1681340463
transform 1 0 -2810 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M62
timestamp 1681340463
transform 1 0 -2352 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M63
timestamp 1681340463
transform -1 0 -1746 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M64
timestamp 1681340463
transform 1 0 -1288 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M65
timestamp 1681340463
transform 1 0 -682 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M66
timestamp 1681340463
transform 1 0 -2810 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M67
timestamp 1681340463
transform 1 0 -2352 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M68
timestamp 1681340463
transform 1 0 -1746 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M69
timestamp 1681340463
transform 1 0 -1288 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M71
timestamp 1681382701
transform 1 0 786 0 1 -3405
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M72
timestamp 1681382701
transform 1 0 1244 0 1 -3405
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M73
timestamp 1681382701
transform 1 0 2914 0 1 -3405
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M74
timestamp 1681382701
transform 1 0 3372 0 1 -3405
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_SMRSPQ  M81
timestamp 1681382701
transform 1 0 172 0 1 -3405
box -108 -557 108 557
use sky130_fd_pr__nfet_01v8_lvt_SMRSPQ  M82
timestamp 1681382701
transform 1 0 330 0 1 -3405
box -108 -557 108 557
use sky130_fd_pr__nfet_01v8_lvt_SMRSPQ  M83
timestamp 1681382701
transform 1 0 2300 0 1 -3405
box -108 -557 108 557
use sky130_fd_pr__nfet_01v8_lvt_SMRSPQ  M84
timestamp 1681382701
transform 1 0 2458 0 1 -3405
box -108 -557 108 557
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M91
timestamp 1681382244
transform 1 0 3214 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M92
timestamp 1681382244
transform 1 0 3672 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M93
timestamp 1681382244
transform 1 0 1086 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M94
timestamp 1681382244
transform 1 0 1544 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M101
timestamp 1681382244
transform 1 0 22 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M102
timestamp 1681382244
transform 1 0 480 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M103
timestamp 1681382244
transform 1 0 2150 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M104
timestamp 1681382244
transform 1 0 2608 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__nfet_01v8_D8YEEC  M111
timestamp 1681382244
transform 1 0 1006 0 1 -4853
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_D8YEEC  M112
timestamp 1681382244
transform 1 0 1612 0 1 -4853
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_D8YEEC  M113
timestamp 1681382244
transform 1 0 2070 0 1 -4853
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_D8YEEC  M114
timestamp 1681382244
transform 1 0 2676 0 1 -4853
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M610
timestamp 1681340463
transform 1 0 -682 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q3 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1671334046
transform 1 0 -3018 0 1 -4856
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q4
timestamp 1671334046
transform 1 0 -1824 0 1 -4856
box 0 0 796 796
<< labels >>
flabel metal1 -5400 -4356 -4896 -2780 0 FreeMono 1280 90 0 0 iin
port 3 nsew
flabel metal2 -5400 -1232 4348 -764 0 FreeMono 1280 0 0 0 vdd
port 0 nsew
flabel metal2 -5400 -5888 4348 -5420 0 FreeMono 1280 0 0 0 vss
port 1 nsew
flabel metal1 4174 -4992 4348 -4192 0 FreeMono 960 90 0 0 vtemp
port 2 nsew
<< end >>
