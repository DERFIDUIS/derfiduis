magic
tech sky130A
timestamp 1680390383
<< pwell >>
rect -133 -205 133 205
<< nmoslvt >>
rect -35 -100 35 100
<< ndiff >>
rect -64 94 -35 100
rect -64 -94 -58 94
rect -41 -94 -35 94
rect -64 -100 -35 -94
rect 35 94 64 100
rect 35 -94 41 94
rect 58 -94 64 94
rect 35 -100 64 -94
<< ndiffc >>
rect -58 -94 -41 94
rect 41 -94 58 94
<< psubdiff >>
rect -115 170 -67 187
rect 67 170 115 187
rect -115 139 -98 170
rect 98 139 115 170
rect -115 -170 -98 -139
rect 98 -170 115 -139
rect -115 -187 -67 -170
rect 67 -187 115 -170
<< psubdiffcont >>
rect -67 170 67 187
rect -115 -139 -98 139
rect 98 -139 115 139
rect -67 -187 67 -170
<< poly >>
rect -35 136 35 144
rect -35 119 -27 136
rect 27 119 35 136
rect -35 100 35 119
rect -35 -119 35 -100
rect -35 -136 -27 -119
rect 27 -136 35 -119
rect -35 -144 35 -136
<< polycont >>
rect -27 119 27 136
rect -27 -136 27 -119
<< locali >>
rect -115 170 -67 187
rect 67 170 115 187
rect -115 139 -98 170
rect 98 139 115 170
rect -35 119 -27 136
rect 27 119 35 136
rect -58 94 -41 102
rect -58 -102 -41 -94
rect 41 94 58 102
rect 41 -102 58 -94
rect -35 -136 -27 -119
rect 27 -136 35 -119
rect -115 -170 -98 -139
rect 98 -170 115 -139
rect -115 -187 -67 -170
rect 67 -187 115 -170
<< viali >>
rect -27 119 27 136
rect -58 -94 -41 94
rect 41 -94 58 94
rect -27 -136 27 -119
<< metal1 >>
rect -33 136 33 139
rect -33 119 -27 136
rect 27 119 33 136
rect -33 116 33 119
rect -61 94 -38 100
rect -61 -94 -58 94
rect -41 -94 -38 94
rect -61 -100 -38 -94
rect 38 94 61 100
rect 38 -94 41 94
rect 58 -94 61 94
rect 38 -100 61 -94
rect -33 -119 33 -116
rect -33 -136 -27 -119
rect 27 -136 33 -119
rect -33 -139 33 -136
<< properties >>
string FIXED_BBOX -106 -178 106 178
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.0 l 0.7 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
