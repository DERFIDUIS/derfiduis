magic
tech sky130A
magscale 1 2
timestamp 1681069304
<< ndiff >>
rect 176 526 178 1526
<< psubdiff >>
rect 112 1472 176 1526
rect 112 1438 116 1472
rect 150 1438 176 1472
rect 112 1404 176 1438
rect 112 1370 116 1404
rect 150 1370 176 1404
rect 112 1336 176 1370
rect 112 1302 116 1336
rect 150 1302 176 1336
rect 112 1268 176 1302
rect 112 1234 116 1268
rect 150 1234 176 1268
rect 112 1200 176 1234
rect 112 1166 116 1200
rect 150 1166 176 1200
rect 112 1132 176 1166
rect 112 1098 116 1132
rect 150 1098 176 1132
rect 112 1064 176 1098
rect 112 1030 116 1064
rect 150 1030 176 1064
rect 112 996 176 1030
rect 112 962 116 996
rect 150 962 176 996
rect 112 928 176 962
rect 112 894 116 928
rect 150 894 176 928
rect 112 860 176 894
rect 112 826 116 860
rect 150 826 176 860
rect 112 792 176 826
rect 112 758 116 792
rect 150 758 176 792
rect 112 724 176 758
rect 112 690 116 724
rect 150 690 176 724
rect 112 656 176 690
rect 112 622 116 656
rect 150 622 176 656
rect 112 588 176 622
rect 112 554 116 588
rect 150 554 176 588
rect 112 526 176 554
<< psubdiffcont >>
rect 116 1438 150 1472
rect 116 1370 150 1404
rect 116 1302 150 1336
rect 116 1234 150 1268
rect 116 1166 150 1200
rect 116 1098 150 1132
rect 116 1030 150 1064
rect 116 962 150 996
rect 116 894 150 928
rect 116 826 150 860
rect 116 758 150 792
rect 116 690 150 724
rect 116 622 150 656
rect 116 554 150 588
<< locali >>
rect 116 1514 150 1530
rect 116 522 150 538
<< viali >>
rect 116 1472 150 1514
rect 116 1438 150 1472
rect 116 1404 150 1438
rect 116 1370 150 1404
rect 116 1336 150 1370
rect 116 1302 150 1336
rect 116 1268 150 1302
rect 116 1234 150 1268
rect 116 1200 150 1234
rect 116 1166 150 1200
rect 116 1132 150 1166
rect 116 1098 150 1132
rect 116 1064 150 1098
rect 116 1030 150 1064
rect 116 996 150 1030
rect 116 962 150 996
rect 116 928 150 962
rect 116 894 150 928
rect 116 860 150 894
rect 116 826 150 860
rect 116 792 150 826
rect 116 758 150 792
rect 116 724 150 758
rect 116 690 150 724
rect 116 656 150 690
rect 116 622 150 656
rect 116 588 150 622
rect 116 554 150 588
rect 116 538 150 554
<< metal1 >>
rect 184 2126 318 2132
rect 184 1684 190 2126
rect 312 1684 318 2126
rect 184 1678 318 1684
rect 224 1558 280 1678
rect -426 1520 42 1526
rect -426 532 -98 1520
rect 36 532 42 1520
rect -426 526 42 532
rect 100 1514 156 1526
rect 388 1520 856 1526
rect 100 538 116 1514
rect 150 538 156 1514
rect 100 396 156 538
rect 184 1514 236 1520
rect 184 532 236 538
rect 266 1514 318 1520
rect 266 532 318 538
rect 388 532 394 1520
rect 528 532 856 1520
rect 388 526 856 532
rect 60 390 194 396
rect 60 -52 66 390
rect 188 -52 194 390
rect 60 -58 194 -52
<< via1 >>
rect 190 1684 312 2126
rect -98 532 36 1520
rect 184 538 236 1514
rect 266 538 318 1514
rect 394 532 528 1520
rect 66 -52 188 390
<< metal2 >>
rect -426 2126 856 2146
rect -426 1684 190 2126
rect 312 1684 856 2126
rect -426 1678 856 1684
rect -104 532 -98 1520
rect 36 1514 236 1520
rect 36 538 184 1514
rect 36 532 236 538
rect 266 1514 394 1520
rect 318 538 394 1514
rect 266 532 394 538
rect 528 532 534 1520
rect -426 390 856 396
rect -426 -52 66 390
rect 188 -52 856 390
rect -426 -72 856 -52
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M1
timestamp 1681062556
transform 1 0 254 0 1 1057
box -76 -557 76 557
<< labels >>
flabel metal1 388 526 856 1526 0 FreeMono 800 0 0 0 outp
port 1 nsew
flabel metal1 -426 526 42 1526 0 FreeMono 800 0 0 0 outn
port 2 nsew
flabel metal2 -426 -72 856 396 0 FreeMono 800 0 0 0 vss
port 0 nsew
flabel metal2 -426 1678 856 2146 0 FreeMono 800 0 0 0 vosc
port 3 nsew
<< end >>
