magic
tech sky130A
magscale 1 2
timestamp 1681251019
<< nwell >>
rect 13884 -3060 13950 -1898
rect 14288 -3060 14402 -1898
rect 14692 -3060 14806 -1898
rect 15096 -3060 15210 -1898
rect 15500 -3060 15614 -1898
rect 15904 -3060 16018 -1898
rect 16356 -3060 16422 -1898
<< ndiff >>
rect 14188 -4436 14190 -3436
rect 14436 -4436 14438 -3436
rect 14524 -4436 14526 -3436
rect 14772 -4436 14774 -3436
rect 14860 -4436 14862 -3436
rect 15108 -4436 15110 -3436
rect 15196 -4436 15198 -3436
rect 15444 -4436 15446 -3436
rect 15532 -4436 15534 -3436
rect 15780 -4436 15782 -3436
rect 15868 -4436 15870 -3436
rect 16116 -4436 16118 -3436
<< pdiff >>
rect 13984 -2960 13986 -1960
rect 14300 -2960 14302 -1960
rect 14388 -2960 14390 -1960
rect 14704 -2960 14706 -1960
rect 14792 -2960 14794 -1960
rect 15108 -2960 15110 -1960
rect 15196 -2960 15198 -1960
rect 15512 -2960 15514 -1960
rect 15600 -2960 15602 -1960
rect 15916 -2960 15918 -1960
rect 16004 -2960 16006 -1960
rect 16320 -2960 16322 -1960
<< psubdiff >>
rect 14124 -3490 14188 -3436
rect 14124 -3524 14128 -3490
rect 14162 -3524 14188 -3490
rect 14124 -3558 14188 -3524
rect 14124 -3592 14128 -3558
rect 14162 -3592 14188 -3558
rect 14124 -3626 14188 -3592
rect 14124 -3660 14128 -3626
rect 14162 -3660 14188 -3626
rect 14124 -3694 14188 -3660
rect 14124 -3728 14128 -3694
rect 14162 -3728 14188 -3694
rect 14124 -3762 14188 -3728
rect 14124 -3796 14128 -3762
rect 14162 -3796 14188 -3762
rect 14124 -3830 14188 -3796
rect 14124 -3864 14128 -3830
rect 14162 -3864 14188 -3830
rect 14124 -3898 14188 -3864
rect 14124 -3932 14128 -3898
rect 14162 -3932 14188 -3898
rect 14124 -3966 14188 -3932
rect 14124 -4000 14128 -3966
rect 14162 -4000 14188 -3966
rect 14124 -4034 14188 -4000
rect 14124 -4068 14128 -4034
rect 14162 -4068 14188 -4034
rect 14124 -4102 14188 -4068
rect 14124 -4136 14128 -4102
rect 14162 -4136 14188 -4102
rect 14124 -4170 14188 -4136
rect 14124 -4204 14128 -4170
rect 14162 -4204 14188 -4170
rect 14124 -4238 14188 -4204
rect 14124 -4272 14128 -4238
rect 14162 -4272 14188 -4238
rect 14124 -4306 14188 -4272
rect 14124 -4340 14128 -4306
rect 14162 -4340 14188 -4306
rect 14124 -4374 14188 -4340
rect 14124 -4408 14128 -4374
rect 14162 -4408 14188 -4374
rect 14124 -4436 14188 -4408
rect 14438 -3464 14524 -3436
rect 14438 -3498 14464 -3464
rect 14498 -3498 14524 -3464
rect 14438 -3532 14524 -3498
rect 14438 -3566 14464 -3532
rect 14498 -3566 14524 -3532
rect 14438 -3600 14524 -3566
rect 14438 -3634 14464 -3600
rect 14498 -3634 14524 -3600
rect 14438 -3668 14524 -3634
rect 14438 -3702 14464 -3668
rect 14498 -3702 14524 -3668
rect 14438 -3736 14524 -3702
rect 14438 -3770 14464 -3736
rect 14498 -3770 14524 -3736
rect 14438 -3804 14524 -3770
rect 14438 -3838 14464 -3804
rect 14498 -3838 14524 -3804
rect 14438 -3872 14524 -3838
rect 14438 -3906 14464 -3872
rect 14498 -3906 14524 -3872
rect 14438 -3940 14524 -3906
rect 14438 -3974 14464 -3940
rect 14498 -3974 14524 -3940
rect 14438 -4008 14524 -3974
rect 14438 -4042 14464 -4008
rect 14498 -4042 14524 -4008
rect 14438 -4076 14524 -4042
rect 14438 -4110 14464 -4076
rect 14498 -4110 14524 -4076
rect 14438 -4144 14524 -4110
rect 14438 -4178 14464 -4144
rect 14498 -4178 14524 -4144
rect 14438 -4212 14524 -4178
rect 14438 -4246 14464 -4212
rect 14498 -4246 14524 -4212
rect 14438 -4280 14524 -4246
rect 14438 -4314 14464 -4280
rect 14498 -4314 14524 -4280
rect 14438 -4348 14524 -4314
rect 14438 -4382 14464 -4348
rect 14498 -4382 14524 -4348
rect 14438 -4436 14524 -4382
rect 14774 -3464 14860 -3436
rect 14774 -3498 14800 -3464
rect 14834 -3498 14860 -3464
rect 14774 -3532 14860 -3498
rect 14774 -3566 14800 -3532
rect 14834 -3566 14860 -3532
rect 14774 -3600 14860 -3566
rect 14774 -3634 14800 -3600
rect 14834 -3634 14860 -3600
rect 14774 -3668 14860 -3634
rect 14774 -3702 14800 -3668
rect 14834 -3702 14860 -3668
rect 14774 -3736 14860 -3702
rect 14774 -3770 14800 -3736
rect 14834 -3770 14860 -3736
rect 14774 -3804 14860 -3770
rect 14774 -3838 14800 -3804
rect 14834 -3838 14860 -3804
rect 14774 -3872 14860 -3838
rect 14774 -3906 14800 -3872
rect 14834 -3906 14860 -3872
rect 14774 -3940 14860 -3906
rect 14774 -3974 14800 -3940
rect 14834 -3974 14860 -3940
rect 14774 -4008 14860 -3974
rect 14774 -4042 14800 -4008
rect 14834 -4042 14860 -4008
rect 14774 -4076 14860 -4042
rect 14774 -4110 14800 -4076
rect 14834 -4110 14860 -4076
rect 14774 -4144 14860 -4110
rect 14774 -4178 14800 -4144
rect 14834 -4178 14860 -4144
rect 14774 -4212 14860 -4178
rect 14774 -4246 14800 -4212
rect 14834 -4246 14860 -4212
rect 14774 -4280 14860 -4246
rect 14774 -4314 14800 -4280
rect 14834 -4314 14860 -4280
rect 14774 -4348 14860 -4314
rect 14774 -4382 14800 -4348
rect 14834 -4382 14860 -4348
rect 14774 -4436 14860 -4382
rect 15110 -3464 15196 -3436
rect 15110 -3498 15136 -3464
rect 15170 -3498 15196 -3464
rect 15110 -3532 15196 -3498
rect 15110 -3566 15136 -3532
rect 15170 -3566 15196 -3532
rect 15110 -3600 15196 -3566
rect 15110 -3634 15136 -3600
rect 15170 -3634 15196 -3600
rect 15110 -3668 15196 -3634
rect 15110 -3702 15136 -3668
rect 15170 -3702 15196 -3668
rect 15110 -3736 15196 -3702
rect 15110 -3770 15136 -3736
rect 15170 -3770 15196 -3736
rect 15110 -3804 15196 -3770
rect 15110 -3838 15136 -3804
rect 15170 -3838 15196 -3804
rect 15110 -3872 15196 -3838
rect 15110 -3906 15136 -3872
rect 15170 -3906 15196 -3872
rect 15110 -3940 15196 -3906
rect 15110 -3974 15136 -3940
rect 15170 -3974 15196 -3940
rect 15110 -4008 15196 -3974
rect 15110 -4042 15136 -4008
rect 15170 -4042 15196 -4008
rect 15110 -4076 15196 -4042
rect 15110 -4110 15136 -4076
rect 15170 -4110 15196 -4076
rect 15110 -4144 15196 -4110
rect 15110 -4178 15136 -4144
rect 15170 -4178 15196 -4144
rect 15110 -4212 15196 -4178
rect 15110 -4246 15136 -4212
rect 15170 -4246 15196 -4212
rect 15110 -4280 15196 -4246
rect 15110 -4314 15136 -4280
rect 15170 -4314 15196 -4280
rect 15110 -4348 15196 -4314
rect 15110 -4382 15136 -4348
rect 15170 -4382 15196 -4348
rect 15110 -4436 15196 -4382
rect 15446 -3464 15532 -3436
rect 15446 -3498 15472 -3464
rect 15506 -3498 15532 -3464
rect 15446 -3532 15532 -3498
rect 15446 -3566 15472 -3532
rect 15506 -3566 15532 -3532
rect 15446 -3600 15532 -3566
rect 15446 -3634 15472 -3600
rect 15506 -3634 15532 -3600
rect 15446 -3668 15532 -3634
rect 15446 -3702 15472 -3668
rect 15506 -3702 15532 -3668
rect 15446 -3736 15532 -3702
rect 15446 -3770 15472 -3736
rect 15506 -3770 15532 -3736
rect 15446 -3804 15532 -3770
rect 15446 -3838 15472 -3804
rect 15506 -3838 15532 -3804
rect 15446 -3872 15532 -3838
rect 15446 -3906 15472 -3872
rect 15506 -3906 15532 -3872
rect 15446 -3940 15532 -3906
rect 15446 -3974 15472 -3940
rect 15506 -3974 15532 -3940
rect 15446 -4008 15532 -3974
rect 15446 -4042 15472 -4008
rect 15506 -4042 15532 -4008
rect 15446 -4076 15532 -4042
rect 15446 -4110 15472 -4076
rect 15506 -4110 15532 -4076
rect 15446 -4144 15532 -4110
rect 15446 -4178 15472 -4144
rect 15506 -4178 15532 -4144
rect 15446 -4212 15532 -4178
rect 15446 -4246 15472 -4212
rect 15506 -4246 15532 -4212
rect 15446 -4280 15532 -4246
rect 15446 -4314 15472 -4280
rect 15506 -4314 15532 -4280
rect 15446 -4348 15532 -4314
rect 15446 -4382 15472 -4348
rect 15506 -4382 15532 -4348
rect 15446 -4436 15532 -4382
rect 15782 -3464 15868 -3436
rect 15782 -3498 15808 -3464
rect 15842 -3498 15868 -3464
rect 15782 -3532 15868 -3498
rect 15782 -3566 15808 -3532
rect 15842 -3566 15868 -3532
rect 15782 -3600 15868 -3566
rect 15782 -3634 15808 -3600
rect 15842 -3634 15868 -3600
rect 15782 -3668 15868 -3634
rect 15782 -3702 15808 -3668
rect 15842 -3702 15868 -3668
rect 15782 -3736 15868 -3702
rect 15782 -3770 15808 -3736
rect 15842 -3770 15868 -3736
rect 15782 -3804 15868 -3770
rect 15782 -3838 15808 -3804
rect 15842 -3838 15868 -3804
rect 15782 -3872 15868 -3838
rect 15782 -3906 15808 -3872
rect 15842 -3906 15868 -3872
rect 15782 -3940 15868 -3906
rect 15782 -3974 15808 -3940
rect 15842 -3974 15868 -3940
rect 15782 -4008 15868 -3974
rect 15782 -4042 15808 -4008
rect 15842 -4042 15868 -4008
rect 15782 -4076 15868 -4042
rect 15782 -4110 15808 -4076
rect 15842 -4110 15868 -4076
rect 15782 -4144 15868 -4110
rect 15782 -4178 15808 -4144
rect 15842 -4178 15868 -4144
rect 15782 -4212 15868 -4178
rect 15782 -4246 15808 -4212
rect 15842 -4246 15868 -4212
rect 15782 -4280 15868 -4246
rect 15782 -4314 15808 -4280
rect 15842 -4314 15868 -4280
rect 15782 -4348 15868 -4314
rect 15782 -4382 15808 -4348
rect 15842 -4382 15868 -4348
rect 15782 -4436 15868 -4382
rect 16118 -3464 16182 -3436
rect 16118 -3498 16144 -3464
rect 16178 -3498 16182 -3464
rect 16118 -3532 16182 -3498
rect 16118 -3566 16144 -3532
rect 16178 -3566 16182 -3532
rect 16118 -3600 16182 -3566
rect 16118 -3634 16144 -3600
rect 16178 -3634 16182 -3600
rect 16118 -3668 16182 -3634
rect 16118 -3702 16144 -3668
rect 16178 -3702 16182 -3668
rect 16118 -3736 16182 -3702
rect 16118 -3770 16144 -3736
rect 16178 -3770 16182 -3736
rect 16118 -3804 16182 -3770
rect 16118 -3838 16144 -3804
rect 16178 -3838 16182 -3804
rect 16118 -3872 16182 -3838
rect 16118 -3906 16144 -3872
rect 16178 -3906 16182 -3872
rect 16118 -3940 16182 -3906
rect 16118 -3974 16144 -3940
rect 16178 -3974 16182 -3940
rect 16118 -4008 16182 -3974
rect 16118 -4042 16144 -4008
rect 16178 -4042 16182 -4008
rect 16118 -4076 16182 -4042
rect 16118 -4110 16144 -4076
rect 16178 -4110 16182 -4076
rect 16118 -4144 16182 -4110
rect 16118 -4178 16144 -4144
rect 16178 -4178 16182 -4144
rect 16118 -4212 16182 -4178
rect 16118 -4246 16144 -4212
rect 16178 -4246 16182 -4212
rect 16118 -4280 16182 -4246
rect 16118 -4314 16144 -4280
rect 16178 -4314 16182 -4280
rect 16118 -4348 16182 -4314
rect 16118 -4382 16144 -4348
rect 16178 -4382 16182 -4348
rect 16118 -4436 16182 -4382
<< nsubdiff >>
rect 13920 -2014 13984 -1960
rect 13920 -2048 13924 -2014
rect 13958 -2048 13984 -2014
rect 13920 -2082 13984 -2048
rect 13920 -2116 13924 -2082
rect 13958 -2116 13984 -2082
rect 13920 -2150 13984 -2116
rect 13920 -2184 13924 -2150
rect 13958 -2184 13984 -2150
rect 13920 -2218 13984 -2184
rect 13920 -2252 13924 -2218
rect 13958 -2252 13984 -2218
rect 13920 -2286 13984 -2252
rect 13920 -2320 13924 -2286
rect 13958 -2320 13984 -2286
rect 13920 -2354 13984 -2320
rect 13920 -2388 13924 -2354
rect 13958 -2388 13984 -2354
rect 13920 -2422 13984 -2388
rect 13920 -2456 13924 -2422
rect 13958 -2456 13984 -2422
rect 13920 -2490 13984 -2456
rect 13920 -2524 13924 -2490
rect 13958 -2524 13984 -2490
rect 13920 -2558 13984 -2524
rect 13920 -2592 13924 -2558
rect 13958 -2592 13984 -2558
rect 13920 -2626 13984 -2592
rect 13920 -2660 13924 -2626
rect 13958 -2660 13984 -2626
rect 13920 -2694 13984 -2660
rect 13920 -2728 13924 -2694
rect 13958 -2728 13984 -2694
rect 13920 -2762 13984 -2728
rect 13920 -2796 13924 -2762
rect 13958 -2796 13984 -2762
rect 13920 -2830 13984 -2796
rect 13920 -2864 13924 -2830
rect 13958 -2864 13984 -2830
rect 13920 -2898 13984 -2864
rect 13920 -2932 13924 -2898
rect 13958 -2932 13984 -2898
rect 13920 -2960 13984 -2932
rect 14302 -1988 14388 -1960
rect 14302 -2022 14328 -1988
rect 14362 -2022 14388 -1988
rect 14302 -2056 14388 -2022
rect 14302 -2090 14328 -2056
rect 14362 -2090 14388 -2056
rect 14302 -2124 14388 -2090
rect 14302 -2158 14328 -2124
rect 14362 -2158 14388 -2124
rect 14302 -2192 14388 -2158
rect 14302 -2226 14328 -2192
rect 14362 -2226 14388 -2192
rect 14302 -2260 14388 -2226
rect 14302 -2294 14328 -2260
rect 14362 -2294 14388 -2260
rect 14302 -2328 14388 -2294
rect 14302 -2362 14328 -2328
rect 14362 -2362 14388 -2328
rect 14302 -2396 14388 -2362
rect 14302 -2430 14328 -2396
rect 14362 -2430 14388 -2396
rect 14302 -2464 14388 -2430
rect 14302 -2498 14328 -2464
rect 14362 -2498 14388 -2464
rect 14302 -2532 14388 -2498
rect 14302 -2566 14328 -2532
rect 14362 -2566 14388 -2532
rect 14302 -2600 14388 -2566
rect 14302 -2634 14328 -2600
rect 14362 -2634 14388 -2600
rect 14302 -2668 14388 -2634
rect 14302 -2702 14328 -2668
rect 14362 -2702 14388 -2668
rect 14302 -2736 14388 -2702
rect 14302 -2770 14328 -2736
rect 14362 -2770 14388 -2736
rect 14302 -2804 14388 -2770
rect 14302 -2838 14328 -2804
rect 14362 -2838 14388 -2804
rect 14302 -2872 14388 -2838
rect 14302 -2906 14328 -2872
rect 14362 -2906 14388 -2872
rect 14302 -2960 14388 -2906
rect 14706 -1988 14792 -1960
rect 14706 -2022 14732 -1988
rect 14766 -2022 14792 -1988
rect 14706 -2056 14792 -2022
rect 14706 -2090 14732 -2056
rect 14766 -2090 14792 -2056
rect 14706 -2124 14792 -2090
rect 14706 -2158 14732 -2124
rect 14766 -2158 14792 -2124
rect 14706 -2192 14792 -2158
rect 14706 -2226 14732 -2192
rect 14766 -2226 14792 -2192
rect 14706 -2260 14792 -2226
rect 14706 -2294 14732 -2260
rect 14766 -2294 14792 -2260
rect 14706 -2328 14792 -2294
rect 14706 -2362 14732 -2328
rect 14766 -2362 14792 -2328
rect 14706 -2396 14792 -2362
rect 14706 -2430 14732 -2396
rect 14766 -2430 14792 -2396
rect 14706 -2464 14792 -2430
rect 14706 -2498 14732 -2464
rect 14766 -2498 14792 -2464
rect 14706 -2532 14792 -2498
rect 14706 -2566 14732 -2532
rect 14766 -2566 14792 -2532
rect 14706 -2600 14792 -2566
rect 14706 -2634 14732 -2600
rect 14766 -2634 14792 -2600
rect 14706 -2668 14792 -2634
rect 14706 -2702 14732 -2668
rect 14766 -2702 14792 -2668
rect 14706 -2736 14792 -2702
rect 14706 -2770 14732 -2736
rect 14766 -2770 14792 -2736
rect 14706 -2804 14792 -2770
rect 14706 -2838 14732 -2804
rect 14766 -2838 14792 -2804
rect 14706 -2872 14792 -2838
rect 14706 -2906 14732 -2872
rect 14766 -2906 14792 -2872
rect 14706 -2960 14792 -2906
rect 15110 -1988 15196 -1960
rect 15110 -2022 15136 -1988
rect 15170 -2022 15196 -1988
rect 15110 -2056 15196 -2022
rect 15110 -2090 15136 -2056
rect 15170 -2090 15196 -2056
rect 15110 -2124 15196 -2090
rect 15110 -2158 15136 -2124
rect 15170 -2158 15196 -2124
rect 15110 -2192 15196 -2158
rect 15110 -2226 15136 -2192
rect 15170 -2226 15196 -2192
rect 15110 -2260 15196 -2226
rect 15110 -2294 15136 -2260
rect 15170 -2294 15196 -2260
rect 15110 -2328 15196 -2294
rect 15110 -2362 15136 -2328
rect 15170 -2362 15196 -2328
rect 15110 -2396 15196 -2362
rect 15110 -2430 15136 -2396
rect 15170 -2430 15196 -2396
rect 15110 -2464 15196 -2430
rect 15110 -2498 15136 -2464
rect 15170 -2498 15196 -2464
rect 15110 -2532 15196 -2498
rect 15110 -2566 15136 -2532
rect 15170 -2566 15196 -2532
rect 15110 -2600 15196 -2566
rect 15110 -2634 15136 -2600
rect 15170 -2634 15196 -2600
rect 15110 -2668 15196 -2634
rect 15110 -2702 15136 -2668
rect 15170 -2702 15196 -2668
rect 15110 -2736 15196 -2702
rect 15110 -2770 15136 -2736
rect 15170 -2770 15196 -2736
rect 15110 -2804 15196 -2770
rect 15110 -2838 15136 -2804
rect 15170 -2838 15196 -2804
rect 15110 -2872 15196 -2838
rect 15110 -2906 15136 -2872
rect 15170 -2906 15196 -2872
rect 15110 -2960 15196 -2906
rect 15514 -1988 15600 -1960
rect 15514 -2022 15540 -1988
rect 15574 -2022 15600 -1988
rect 15514 -2056 15600 -2022
rect 15514 -2090 15540 -2056
rect 15574 -2090 15600 -2056
rect 15514 -2124 15600 -2090
rect 15514 -2158 15540 -2124
rect 15574 -2158 15600 -2124
rect 15514 -2192 15600 -2158
rect 15514 -2226 15540 -2192
rect 15574 -2226 15600 -2192
rect 15514 -2260 15600 -2226
rect 15514 -2294 15540 -2260
rect 15574 -2294 15600 -2260
rect 15514 -2328 15600 -2294
rect 15514 -2362 15540 -2328
rect 15574 -2362 15600 -2328
rect 15514 -2396 15600 -2362
rect 15514 -2430 15540 -2396
rect 15574 -2430 15600 -2396
rect 15514 -2464 15600 -2430
rect 15514 -2498 15540 -2464
rect 15574 -2498 15600 -2464
rect 15514 -2532 15600 -2498
rect 15514 -2566 15540 -2532
rect 15574 -2566 15600 -2532
rect 15514 -2600 15600 -2566
rect 15514 -2634 15540 -2600
rect 15574 -2634 15600 -2600
rect 15514 -2668 15600 -2634
rect 15514 -2702 15540 -2668
rect 15574 -2702 15600 -2668
rect 15514 -2736 15600 -2702
rect 15514 -2770 15540 -2736
rect 15574 -2770 15600 -2736
rect 15514 -2804 15600 -2770
rect 15514 -2838 15540 -2804
rect 15574 -2838 15600 -2804
rect 15514 -2872 15600 -2838
rect 15514 -2906 15540 -2872
rect 15574 -2906 15600 -2872
rect 15514 -2960 15600 -2906
rect 15918 -1988 16004 -1960
rect 15918 -2022 15944 -1988
rect 15978 -2022 16004 -1988
rect 15918 -2056 16004 -2022
rect 15918 -2090 15944 -2056
rect 15978 -2090 16004 -2056
rect 15918 -2124 16004 -2090
rect 15918 -2158 15944 -2124
rect 15978 -2158 16004 -2124
rect 15918 -2192 16004 -2158
rect 15918 -2226 15944 -2192
rect 15978 -2226 16004 -2192
rect 15918 -2260 16004 -2226
rect 15918 -2294 15944 -2260
rect 15978 -2294 16004 -2260
rect 15918 -2328 16004 -2294
rect 15918 -2362 15944 -2328
rect 15978 -2362 16004 -2328
rect 15918 -2396 16004 -2362
rect 15918 -2430 15944 -2396
rect 15978 -2430 16004 -2396
rect 15918 -2464 16004 -2430
rect 15918 -2498 15944 -2464
rect 15978 -2498 16004 -2464
rect 15918 -2532 16004 -2498
rect 15918 -2566 15944 -2532
rect 15978 -2566 16004 -2532
rect 15918 -2600 16004 -2566
rect 15918 -2634 15944 -2600
rect 15978 -2634 16004 -2600
rect 15918 -2668 16004 -2634
rect 15918 -2702 15944 -2668
rect 15978 -2702 16004 -2668
rect 15918 -2736 16004 -2702
rect 15918 -2770 15944 -2736
rect 15978 -2770 16004 -2736
rect 15918 -2804 16004 -2770
rect 15918 -2838 15944 -2804
rect 15978 -2838 16004 -2804
rect 15918 -2872 16004 -2838
rect 15918 -2906 15944 -2872
rect 15978 -2906 16004 -2872
rect 15918 -2960 16004 -2906
rect 16322 -1988 16386 -1960
rect 16322 -2022 16348 -1988
rect 16382 -2022 16386 -1988
rect 16322 -2056 16386 -2022
rect 16322 -2090 16348 -2056
rect 16382 -2090 16386 -2056
rect 16322 -2124 16386 -2090
rect 16322 -2158 16348 -2124
rect 16382 -2158 16386 -2124
rect 16322 -2192 16386 -2158
rect 16322 -2226 16348 -2192
rect 16382 -2226 16386 -2192
rect 16322 -2260 16386 -2226
rect 16322 -2294 16348 -2260
rect 16382 -2294 16386 -2260
rect 16322 -2328 16386 -2294
rect 16322 -2362 16348 -2328
rect 16382 -2362 16386 -2328
rect 16322 -2396 16386 -2362
rect 16322 -2430 16348 -2396
rect 16382 -2430 16386 -2396
rect 16322 -2464 16386 -2430
rect 16322 -2498 16348 -2464
rect 16382 -2498 16386 -2464
rect 16322 -2532 16386 -2498
rect 16322 -2566 16348 -2532
rect 16382 -2566 16386 -2532
rect 16322 -2600 16386 -2566
rect 16322 -2634 16348 -2600
rect 16382 -2634 16386 -2600
rect 16322 -2668 16386 -2634
rect 16322 -2702 16348 -2668
rect 16382 -2702 16386 -2668
rect 16322 -2736 16386 -2702
rect 16322 -2770 16348 -2736
rect 16382 -2770 16386 -2736
rect 16322 -2804 16386 -2770
rect 16322 -2838 16348 -2804
rect 16382 -2838 16386 -2804
rect 16322 -2872 16386 -2838
rect 16322 -2906 16348 -2872
rect 16382 -2906 16386 -2872
rect 16322 -2960 16386 -2906
<< psubdiffcont >>
rect 14128 -3524 14162 -3490
rect 14128 -3592 14162 -3558
rect 14128 -3660 14162 -3626
rect 14128 -3728 14162 -3694
rect 14128 -3796 14162 -3762
rect 14128 -3864 14162 -3830
rect 14128 -3932 14162 -3898
rect 14128 -4000 14162 -3966
rect 14128 -4068 14162 -4034
rect 14128 -4136 14162 -4102
rect 14128 -4204 14162 -4170
rect 14128 -4272 14162 -4238
rect 14128 -4340 14162 -4306
rect 14128 -4408 14162 -4374
rect 14464 -3498 14498 -3464
rect 14464 -3566 14498 -3532
rect 14464 -3634 14498 -3600
rect 14464 -3702 14498 -3668
rect 14464 -3770 14498 -3736
rect 14464 -3838 14498 -3804
rect 14464 -3906 14498 -3872
rect 14464 -3974 14498 -3940
rect 14464 -4042 14498 -4008
rect 14464 -4110 14498 -4076
rect 14464 -4178 14498 -4144
rect 14464 -4246 14498 -4212
rect 14464 -4314 14498 -4280
rect 14464 -4382 14498 -4348
rect 14800 -3498 14834 -3464
rect 14800 -3566 14834 -3532
rect 14800 -3634 14834 -3600
rect 14800 -3702 14834 -3668
rect 14800 -3770 14834 -3736
rect 14800 -3838 14834 -3804
rect 14800 -3906 14834 -3872
rect 14800 -3974 14834 -3940
rect 14800 -4042 14834 -4008
rect 14800 -4110 14834 -4076
rect 14800 -4178 14834 -4144
rect 14800 -4246 14834 -4212
rect 14800 -4314 14834 -4280
rect 14800 -4382 14834 -4348
rect 15136 -3498 15170 -3464
rect 15136 -3566 15170 -3532
rect 15136 -3634 15170 -3600
rect 15136 -3702 15170 -3668
rect 15136 -3770 15170 -3736
rect 15136 -3838 15170 -3804
rect 15136 -3906 15170 -3872
rect 15136 -3974 15170 -3940
rect 15136 -4042 15170 -4008
rect 15136 -4110 15170 -4076
rect 15136 -4178 15170 -4144
rect 15136 -4246 15170 -4212
rect 15136 -4314 15170 -4280
rect 15136 -4382 15170 -4348
rect 15472 -3498 15506 -3464
rect 15472 -3566 15506 -3532
rect 15472 -3634 15506 -3600
rect 15472 -3702 15506 -3668
rect 15472 -3770 15506 -3736
rect 15472 -3838 15506 -3804
rect 15472 -3906 15506 -3872
rect 15472 -3974 15506 -3940
rect 15472 -4042 15506 -4008
rect 15472 -4110 15506 -4076
rect 15472 -4178 15506 -4144
rect 15472 -4246 15506 -4212
rect 15472 -4314 15506 -4280
rect 15472 -4382 15506 -4348
rect 15808 -3498 15842 -3464
rect 15808 -3566 15842 -3532
rect 15808 -3634 15842 -3600
rect 15808 -3702 15842 -3668
rect 15808 -3770 15842 -3736
rect 15808 -3838 15842 -3804
rect 15808 -3906 15842 -3872
rect 15808 -3974 15842 -3940
rect 15808 -4042 15842 -4008
rect 15808 -4110 15842 -4076
rect 15808 -4178 15842 -4144
rect 15808 -4246 15842 -4212
rect 15808 -4314 15842 -4280
rect 15808 -4382 15842 -4348
rect 16144 -3498 16178 -3464
rect 16144 -3566 16178 -3532
rect 16144 -3634 16178 -3600
rect 16144 -3702 16178 -3668
rect 16144 -3770 16178 -3736
rect 16144 -3838 16178 -3804
rect 16144 -3906 16178 -3872
rect 16144 -3974 16178 -3940
rect 16144 -4042 16178 -4008
rect 16144 -4110 16178 -4076
rect 16144 -4178 16178 -4144
rect 16144 -4246 16178 -4212
rect 16144 -4314 16178 -4280
rect 16144 -4382 16178 -4348
<< nsubdiffcont >>
rect 13924 -2048 13958 -2014
rect 13924 -2116 13958 -2082
rect 13924 -2184 13958 -2150
rect 13924 -2252 13958 -2218
rect 13924 -2320 13958 -2286
rect 13924 -2388 13958 -2354
rect 13924 -2456 13958 -2422
rect 13924 -2524 13958 -2490
rect 13924 -2592 13958 -2558
rect 13924 -2660 13958 -2626
rect 13924 -2728 13958 -2694
rect 13924 -2796 13958 -2762
rect 13924 -2864 13958 -2830
rect 13924 -2932 13958 -2898
rect 14328 -2022 14362 -1988
rect 14328 -2090 14362 -2056
rect 14328 -2158 14362 -2124
rect 14328 -2226 14362 -2192
rect 14328 -2294 14362 -2260
rect 14328 -2362 14362 -2328
rect 14328 -2430 14362 -2396
rect 14328 -2498 14362 -2464
rect 14328 -2566 14362 -2532
rect 14328 -2634 14362 -2600
rect 14328 -2702 14362 -2668
rect 14328 -2770 14362 -2736
rect 14328 -2838 14362 -2804
rect 14328 -2906 14362 -2872
rect 14732 -2022 14766 -1988
rect 14732 -2090 14766 -2056
rect 14732 -2158 14766 -2124
rect 14732 -2226 14766 -2192
rect 14732 -2294 14766 -2260
rect 14732 -2362 14766 -2328
rect 14732 -2430 14766 -2396
rect 14732 -2498 14766 -2464
rect 14732 -2566 14766 -2532
rect 14732 -2634 14766 -2600
rect 14732 -2702 14766 -2668
rect 14732 -2770 14766 -2736
rect 14732 -2838 14766 -2804
rect 14732 -2906 14766 -2872
rect 15136 -2022 15170 -1988
rect 15136 -2090 15170 -2056
rect 15136 -2158 15170 -2124
rect 15136 -2226 15170 -2192
rect 15136 -2294 15170 -2260
rect 15136 -2362 15170 -2328
rect 15136 -2430 15170 -2396
rect 15136 -2498 15170 -2464
rect 15136 -2566 15170 -2532
rect 15136 -2634 15170 -2600
rect 15136 -2702 15170 -2668
rect 15136 -2770 15170 -2736
rect 15136 -2838 15170 -2804
rect 15136 -2906 15170 -2872
rect 15540 -2022 15574 -1988
rect 15540 -2090 15574 -2056
rect 15540 -2158 15574 -2124
rect 15540 -2226 15574 -2192
rect 15540 -2294 15574 -2260
rect 15540 -2362 15574 -2328
rect 15540 -2430 15574 -2396
rect 15540 -2498 15574 -2464
rect 15540 -2566 15574 -2532
rect 15540 -2634 15574 -2600
rect 15540 -2702 15574 -2668
rect 15540 -2770 15574 -2736
rect 15540 -2838 15574 -2804
rect 15540 -2906 15574 -2872
rect 15944 -2022 15978 -1988
rect 15944 -2090 15978 -2056
rect 15944 -2158 15978 -2124
rect 15944 -2226 15978 -2192
rect 15944 -2294 15978 -2260
rect 15944 -2362 15978 -2328
rect 15944 -2430 15978 -2396
rect 15944 -2498 15978 -2464
rect 15944 -2566 15978 -2532
rect 15944 -2634 15978 -2600
rect 15944 -2702 15978 -2668
rect 15944 -2770 15978 -2736
rect 15944 -2838 15978 -2804
rect 15944 -2906 15978 -2872
rect 16348 -2022 16382 -1988
rect 16348 -2090 16382 -2056
rect 16348 -2158 16382 -2124
rect 16348 -2226 16382 -2192
rect 16348 -2294 16382 -2260
rect 16348 -2362 16382 -2328
rect 16348 -2430 16382 -2396
rect 16348 -2498 16382 -2464
rect 16348 -2566 16382 -2532
rect 16348 -2634 16382 -2600
rect 16348 -2702 16382 -2668
rect 16348 -2770 16382 -2736
rect 16348 -2838 16382 -2804
rect 16348 -2906 16382 -2872
<< poly >>
rect 14298 -3414 14328 -3348
rect 14634 -3414 14664 -3348
rect 14970 -3414 15000 -3348
rect 15306 -3414 15336 -3348
rect 15642 -3414 15672 -3348
rect 15978 -3414 16008 -3348
<< locali >>
rect 13924 -1972 13958 -1956
rect 13924 -2964 13958 -2948
rect 14328 -1972 14362 -1956
rect 14328 -2964 14362 -2948
rect 14732 -1972 14766 -1956
rect 14732 -2964 14766 -2948
rect 15136 -1972 15170 -1956
rect 15136 -2964 15170 -2948
rect 15540 -1972 15574 -1956
rect 15540 -2964 15574 -2948
rect 15944 -1972 15978 -1956
rect 15944 -2964 15978 -2948
rect 16348 -1972 16382 -1956
rect 16348 -2964 16382 -2948
rect 14298 -3398 14328 -3364
rect 14634 -3398 14664 -3364
rect 14970 -3398 15000 -3364
rect 15306 -3398 15336 -3364
rect 15642 -3398 15672 -3364
rect 15978 -3398 16008 -3364
rect 14128 -3490 14162 -3432
rect 14128 -3558 14162 -3524
rect 14128 -3626 14162 -3592
rect 14128 -3694 14162 -3660
rect 14128 -3736 14162 -3728
rect 14128 -4440 14162 -4424
rect 14464 -3464 14498 -3432
rect 14464 -3532 14498 -3498
rect 14464 -3600 14498 -3566
rect 14464 -3668 14498 -3634
rect 14464 -3736 14498 -3702
rect 14464 -4440 14498 -4424
rect 14800 -3464 14834 -3432
rect 14800 -3532 14834 -3498
rect 14800 -3600 14834 -3566
rect 14800 -3668 14834 -3634
rect 14800 -3736 14834 -3702
rect 14800 -4440 14834 -4424
rect 15136 -3464 15170 -3432
rect 15136 -3532 15170 -3498
rect 15136 -3600 15170 -3566
rect 15136 -3668 15170 -3634
rect 15136 -3736 15170 -3702
rect 15136 -4440 15170 -4424
rect 15472 -3464 15506 -3432
rect 15472 -3532 15506 -3498
rect 15472 -3600 15506 -3566
rect 15472 -3668 15506 -3634
rect 15472 -3736 15506 -3702
rect 15472 -4440 15506 -4424
rect 15808 -3464 15842 -3432
rect 15808 -3532 15842 -3498
rect 15808 -3600 15842 -3566
rect 15808 -3668 15842 -3634
rect 15808 -3736 15842 -3702
rect 15808 -4440 15842 -4424
rect 16144 -3464 16178 -3432
rect 16144 -3532 16178 -3498
rect 16144 -3600 16178 -3566
rect 16144 -3668 16178 -3634
rect 16144 -3736 16178 -3702
rect 16144 -4440 16178 -4424
<< viali >>
rect 13924 -2014 13958 -1972
rect 13924 -2048 13958 -2014
rect 13924 -2082 13958 -2048
rect 13924 -2116 13958 -2082
rect 13924 -2150 13958 -2116
rect 13924 -2184 13958 -2150
rect 13924 -2218 13958 -2184
rect 13924 -2252 13958 -2218
rect 13924 -2286 13958 -2252
rect 13924 -2320 13958 -2286
rect 13924 -2354 13958 -2320
rect 13924 -2388 13958 -2354
rect 13924 -2422 13958 -2388
rect 13924 -2456 13958 -2422
rect 13924 -2490 13958 -2456
rect 13924 -2524 13958 -2490
rect 13924 -2558 13958 -2524
rect 13924 -2592 13958 -2558
rect 13924 -2626 13958 -2592
rect 13924 -2660 13958 -2626
rect 13924 -2694 13958 -2660
rect 13924 -2728 13958 -2694
rect 13924 -2762 13958 -2728
rect 13924 -2796 13958 -2762
rect 13924 -2830 13958 -2796
rect 13924 -2864 13958 -2830
rect 13924 -2898 13958 -2864
rect 13924 -2932 13958 -2898
rect 13924 -2948 13958 -2932
rect 14328 -1988 14362 -1972
rect 14328 -2022 14362 -1988
rect 14328 -2056 14362 -2022
rect 14328 -2090 14362 -2056
rect 14328 -2124 14362 -2090
rect 14328 -2158 14362 -2124
rect 14328 -2192 14362 -2158
rect 14328 -2226 14362 -2192
rect 14328 -2260 14362 -2226
rect 14328 -2294 14362 -2260
rect 14328 -2328 14362 -2294
rect 14328 -2362 14362 -2328
rect 14328 -2396 14362 -2362
rect 14328 -2430 14362 -2396
rect 14328 -2464 14362 -2430
rect 14328 -2498 14362 -2464
rect 14328 -2532 14362 -2498
rect 14328 -2566 14362 -2532
rect 14328 -2600 14362 -2566
rect 14328 -2634 14362 -2600
rect 14328 -2668 14362 -2634
rect 14328 -2702 14362 -2668
rect 14328 -2736 14362 -2702
rect 14328 -2770 14362 -2736
rect 14328 -2804 14362 -2770
rect 14328 -2838 14362 -2804
rect 14328 -2872 14362 -2838
rect 14328 -2906 14362 -2872
rect 14328 -2948 14362 -2906
rect 14732 -1988 14766 -1972
rect 14732 -2022 14766 -1988
rect 14732 -2056 14766 -2022
rect 14732 -2090 14766 -2056
rect 14732 -2124 14766 -2090
rect 14732 -2158 14766 -2124
rect 14732 -2192 14766 -2158
rect 14732 -2226 14766 -2192
rect 14732 -2260 14766 -2226
rect 14732 -2294 14766 -2260
rect 14732 -2328 14766 -2294
rect 14732 -2362 14766 -2328
rect 14732 -2396 14766 -2362
rect 14732 -2430 14766 -2396
rect 14732 -2464 14766 -2430
rect 14732 -2498 14766 -2464
rect 14732 -2532 14766 -2498
rect 14732 -2566 14766 -2532
rect 14732 -2600 14766 -2566
rect 14732 -2634 14766 -2600
rect 14732 -2668 14766 -2634
rect 14732 -2702 14766 -2668
rect 14732 -2736 14766 -2702
rect 14732 -2770 14766 -2736
rect 14732 -2804 14766 -2770
rect 14732 -2838 14766 -2804
rect 14732 -2872 14766 -2838
rect 14732 -2906 14766 -2872
rect 14732 -2948 14766 -2906
rect 15136 -1988 15170 -1972
rect 15136 -2022 15170 -1988
rect 15136 -2056 15170 -2022
rect 15136 -2090 15170 -2056
rect 15136 -2124 15170 -2090
rect 15136 -2158 15170 -2124
rect 15136 -2192 15170 -2158
rect 15136 -2226 15170 -2192
rect 15136 -2260 15170 -2226
rect 15136 -2294 15170 -2260
rect 15136 -2328 15170 -2294
rect 15136 -2362 15170 -2328
rect 15136 -2396 15170 -2362
rect 15136 -2430 15170 -2396
rect 15136 -2464 15170 -2430
rect 15136 -2498 15170 -2464
rect 15136 -2532 15170 -2498
rect 15136 -2566 15170 -2532
rect 15136 -2600 15170 -2566
rect 15136 -2634 15170 -2600
rect 15136 -2668 15170 -2634
rect 15136 -2702 15170 -2668
rect 15136 -2736 15170 -2702
rect 15136 -2770 15170 -2736
rect 15136 -2804 15170 -2770
rect 15136 -2838 15170 -2804
rect 15136 -2872 15170 -2838
rect 15136 -2906 15170 -2872
rect 15136 -2948 15170 -2906
rect 15540 -1988 15574 -1972
rect 15540 -2022 15574 -1988
rect 15540 -2056 15574 -2022
rect 15540 -2090 15574 -2056
rect 15540 -2124 15574 -2090
rect 15540 -2158 15574 -2124
rect 15540 -2192 15574 -2158
rect 15540 -2226 15574 -2192
rect 15540 -2260 15574 -2226
rect 15540 -2294 15574 -2260
rect 15540 -2328 15574 -2294
rect 15540 -2362 15574 -2328
rect 15540 -2396 15574 -2362
rect 15540 -2430 15574 -2396
rect 15540 -2464 15574 -2430
rect 15540 -2498 15574 -2464
rect 15540 -2532 15574 -2498
rect 15540 -2566 15574 -2532
rect 15540 -2600 15574 -2566
rect 15540 -2634 15574 -2600
rect 15540 -2668 15574 -2634
rect 15540 -2702 15574 -2668
rect 15540 -2736 15574 -2702
rect 15540 -2770 15574 -2736
rect 15540 -2804 15574 -2770
rect 15540 -2838 15574 -2804
rect 15540 -2872 15574 -2838
rect 15540 -2906 15574 -2872
rect 15540 -2948 15574 -2906
rect 15944 -1988 15978 -1972
rect 15944 -2022 15978 -1988
rect 15944 -2056 15978 -2022
rect 15944 -2090 15978 -2056
rect 15944 -2124 15978 -2090
rect 15944 -2158 15978 -2124
rect 15944 -2192 15978 -2158
rect 15944 -2226 15978 -2192
rect 15944 -2260 15978 -2226
rect 15944 -2294 15978 -2260
rect 15944 -2328 15978 -2294
rect 15944 -2362 15978 -2328
rect 15944 -2396 15978 -2362
rect 15944 -2430 15978 -2396
rect 15944 -2464 15978 -2430
rect 15944 -2498 15978 -2464
rect 15944 -2532 15978 -2498
rect 15944 -2566 15978 -2532
rect 15944 -2600 15978 -2566
rect 15944 -2634 15978 -2600
rect 15944 -2668 15978 -2634
rect 15944 -2702 15978 -2668
rect 15944 -2736 15978 -2702
rect 15944 -2770 15978 -2736
rect 15944 -2804 15978 -2770
rect 15944 -2838 15978 -2804
rect 15944 -2872 15978 -2838
rect 15944 -2906 15978 -2872
rect 15944 -2948 15978 -2906
rect 16348 -1988 16382 -1972
rect 16348 -2022 16382 -1988
rect 16348 -2056 16382 -2022
rect 16348 -2090 16382 -2056
rect 16348 -2124 16382 -2090
rect 16348 -2158 16382 -2124
rect 16348 -2192 16382 -2158
rect 16348 -2226 16382 -2192
rect 16348 -2260 16382 -2226
rect 16348 -2294 16382 -2260
rect 16348 -2328 16382 -2294
rect 16348 -2362 16382 -2328
rect 16348 -2396 16382 -2362
rect 16348 -2430 16382 -2396
rect 16348 -2464 16382 -2430
rect 16348 -2498 16382 -2464
rect 16348 -2532 16382 -2498
rect 16348 -2566 16382 -2532
rect 16348 -2600 16382 -2566
rect 16348 -2634 16382 -2600
rect 16348 -2668 16382 -2634
rect 16348 -2702 16382 -2668
rect 16348 -2736 16382 -2702
rect 16348 -2770 16382 -2736
rect 16348 -2804 16382 -2770
rect 16348 -2838 16382 -2804
rect 16348 -2872 16382 -2838
rect 16348 -2906 16382 -2872
rect 16348 -2948 16382 -2906
rect 14128 -3762 14162 -3736
rect 14128 -3796 14162 -3762
rect 14128 -3830 14162 -3796
rect 14128 -3864 14162 -3830
rect 14128 -3898 14162 -3864
rect 14128 -3932 14162 -3898
rect 14128 -3966 14162 -3932
rect 14128 -4000 14162 -3966
rect 14128 -4034 14162 -4000
rect 14128 -4068 14162 -4034
rect 14128 -4102 14162 -4068
rect 14128 -4136 14162 -4102
rect 14128 -4170 14162 -4136
rect 14128 -4204 14162 -4170
rect 14128 -4238 14162 -4204
rect 14128 -4272 14162 -4238
rect 14128 -4306 14162 -4272
rect 14128 -4340 14162 -4306
rect 14128 -4374 14162 -4340
rect 14128 -4408 14162 -4374
rect 14128 -4424 14162 -4408
rect 14464 -3770 14498 -3736
rect 14464 -3804 14498 -3770
rect 14464 -3838 14498 -3804
rect 14464 -3872 14498 -3838
rect 14464 -3906 14498 -3872
rect 14464 -3940 14498 -3906
rect 14464 -3974 14498 -3940
rect 14464 -4008 14498 -3974
rect 14464 -4042 14498 -4008
rect 14464 -4076 14498 -4042
rect 14464 -4110 14498 -4076
rect 14464 -4144 14498 -4110
rect 14464 -4178 14498 -4144
rect 14464 -4212 14498 -4178
rect 14464 -4246 14498 -4212
rect 14464 -4280 14498 -4246
rect 14464 -4314 14498 -4280
rect 14464 -4348 14498 -4314
rect 14464 -4382 14498 -4348
rect 14464 -4424 14498 -4382
rect 14800 -3770 14834 -3736
rect 14800 -3804 14834 -3770
rect 14800 -3838 14834 -3804
rect 14800 -3872 14834 -3838
rect 14800 -3906 14834 -3872
rect 14800 -3940 14834 -3906
rect 14800 -3974 14834 -3940
rect 14800 -4008 14834 -3974
rect 14800 -4042 14834 -4008
rect 14800 -4076 14834 -4042
rect 14800 -4110 14834 -4076
rect 14800 -4144 14834 -4110
rect 14800 -4178 14834 -4144
rect 14800 -4212 14834 -4178
rect 14800 -4246 14834 -4212
rect 14800 -4280 14834 -4246
rect 14800 -4314 14834 -4280
rect 14800 -4348 14834 -4314
rect 14800 -4382 14834 -4348
rect 14800 -4424 14834 -4382
rect 15136 -3770 15170 -3736
rect 15136 -3804 15170 -3770
rect 15136 -3838 15170 -3804
rect 15136 -3872 15170 -3838
rect 15136 -3906 15170 -3872
rect 15136 -3940 15170 -3906
rect 15136 -3974 15170 -3940
rect 15136 -4008 15170 -3974
rect 15136 -4042 15170 -4008
rect 15136 -4076 15170 -4042
rect 15136 -4110 15170 -4076
rect 15136 -4144 15170 -4110
rect 15136 -4178 15170 -4144
rect 15136 -4212 15170 -4178
rect 15136 -4246 15170 -4212
rect 15136 -4280 15170 -4246
rect 15136 -4314 15170 -4280
rect 15136 -4348 15170 -4314
rect 15136 -4382 15170 -4348
rect 15136 -4424 15170 -4382
rect 15472 -3770 15506 -3736
rect 15472 -3804 15506 -3770
rect 15472 -3838 15506 -3804
rect 15472 -3872 15506 -3838
rect 15472 -3906 15506 -3872
rect 15472 -3940 15506 -3906
rect 15472 -3974 15506 -3940
rect 15472 -4008 15506 -3974
rect 15472 -4042 15506 -4008
rect 15472 -4076 15506 -4042
rect 15472 -4110 15506 -4076
rect 15472 -4144 15506 -4110
rect 15472 -4178 15506 -4144
rect 15472 -4212 15506 -4178
rect 15472 -4246 15506 -4212
rect 15472 -4280 15506 -4246
rect 15472 -4314 15506 -4280
rect 15472 -4348 15506 -4314
rect 15472 -4382 15506 -4348
rect 15472 -4424 15506 -4382
rect 15808 -3770 15842 -3736
rect 15808 -3804 15842 -3770
rect 15808 -3838 15842 -3804
rect 15808 -3872 15842 -3838
rect 15808 -3906 15842 -3872
rect 15808 -3940 15842 -3906
rect 15808 -3974 15842 -3940
rect 15808 -4008 15842 -3974
rect 15808 -4042 15842 -4008
rect 15808 -4076 15842 -4042
rect 15808 -4110 15842 -4076
rect 15808 -4144 15842 -4110
rect 15808 -4178 15842 -4144
rect 15808 -4212 15842 -4178
rect 15808 -4246 15842 -4212
rect 15808 -4280 15842 -4246
rect 15808 -4314 15842 -4280
rect 15808 -4348 15842 -4314
rect 15808 -4382 15842 -4348
rect 15808 -4424 15842 -4382
rect 16144 -3770 16178 -3736
rect 16144 -3804 16178 -3770
rect 16144 -3838 16178 -3804
rect 16144 -3872 16178 -3838
rect 16144 -3906 16178 -3872
rect 16144 -3940 16178 -3906
rect 16144 -3974 16178 -3940
rect 16144 -4008 16178 -3974
rect 16144 -4042 16178 -4008
rect 16144 -4076 16178 -4042
rect 16144 -4110 16178 -4076
rect 16144 -4144 16178 -4110
rect 16144 -4178 16178 -4144
rect 16144 -4212 16178 -4178
rect 16144 -4246 16178 -4212
rect 16144 -4280 16178 -4246
rect 16144 -4314 16178 -4280
rect 16144 -4348 16178 -4314
rect 16144 -4382 16178 -4348
rect 16144 -4424 16178 -4382
<< metal1 >>
rect 13764 -1498 13876 -1488
rect 13764 -1666 13794 -1498
rect 13850 -1666 13876 -1498
rect 13764 -3248 13876 -1666
rect 13904 -1768 16400 -1762
rect 13904 -1820 13924 -1768
rect 16380 -1820 16400 -1768
rect 13904 -1826 16400 -1820
rect 13904 -1972 14016 -1826
rect 13904 -2948 13924 -1972
rect 13958 -2948 14016 -1972
rect 13904 -2960 14016 -2948
rect 14114 -1972 14172 -1962
rect 14114 -2954 14172 -2948
rect 14288 -1972 14400 -1826
rect 14288 -2948 14328 -1972
rect 14362 -2948 14400 -1972
rect 14288 -2960 14400 -2948
rect 14518 -1972 14576 -1962
rect 14518 -2954 14576 -2948
rect 14692 -1972 14804 -1826
rect 14692 -2948 14732 -1972
rect 14766 -2948 14804 -1972
rect 14692 -2960 14804 -2948
rect 14922 -1972 14980 -1962
rect 14922 -2954 14980 -2948
rect 15096 -1972 15208 -1826
rect 15096 -2948 15136 -1972
rect 15170 -2948 15208 -1972
rect 15096 -2960 15208 -2948
rect 15326 -1972 15384 -1962
rect 15326 -2954 15384 -2948
rect 15500 -1972 15612 -1826
rect 15500 -2948 15540 -1972
rect 15574 -2948 15612 -1972
rect 15500 -2960 15612 -2948
rect 15730 -1972 15788 -1962
rect 15730 -2954 15788 -2948
rect 15904 -1972 16016 -1826
rect 15904 -2948 15944 -1972
rect 15978 -2948 16016 -1972
rect 15904 -2960 16016 -2948
rect 16134 -1972 16192 -1962
rect 16134 -2954 16192 -2948
rect 16288 -1972 16400 -1826
rect 16288 -2948 16348 -1972
rect 16382 -2948 16400 -1972
rect 16288 -2960 16400 -2948
rect 14046 -3060 14240 -3000
rect 14450 -3060 14644 -3000
rect 14118 -3102 14240 -3060
rect 14118 -3108 14368 -3102
rect 14342 -3160 14368 -3108
rect 14118 -3166 14368 -3160
rect 13764 -3306 13876 -3300
rect 14234 -3348 14368 -3166
rect 14480 -3242 14614 -3060
rect 14854 -3102 15048 -3000
rect 14854 -3108 15078 -3102
rect 14854 -3166 15078 -3160
rect 14480 -3248 14728 -3242
rect 14704 -3300 14728 -3248
rect 14480 -3306 14728 -3300
rect 14234 -3404 14392 -3348
rect 14570 -3404 14728 -3306
rect 14906 -3404 15064 -3166
rect 15258 -3242 15452 -3000
rect 15662 -3102 15856 -3000
rect 15608 -3108 15856 -3102
rect 15832 -3160 15856 -3108
rect 15608 -3166 15856 -3160
rect 16066 -3078 16260 -3000
rect 15234 -3248 15458 -3242
rect 15234 -3306 15458 -3300
rect 15242 -3404 15400 -3306
rect 15608 -3348 15720 -3166
rect 16066 -3242 16186 -3078
rect 15954 -3248 16186 -3242
rect 16178 -3300 16186 -3248
rect 15954 -3306 16186 -3300
rect 16294 -3108 16406 -3102
rect 15954 -3348 16072 -3306
rect 15578 -3404 15736 -3348
rect 15914 -3404 16072 -3348
rect 8712 -3756 9216 -3706
rect 8712 -4046 9086 -3756
rect 9198 -4046 9216 -3756
rect 8712 -4564 9216 -4046
rect 14106 -3728 14162 -3436
rect 14190 -3442 14248 -3436
rect 14190 -3706 14248 -3700
rect 14378 -3442 14436 -3436
rect 14378 -3706 14436 -3700
rect 14106 -3736 14168 -3728
rect 14464 -3730 14498 -3436
rect 14526 -3442 14584 -3436
rect 14526 -3706 14584 -3700
rect 14714 -3442 14772 -3436
rect 14714 -3706 14772 -3700
rect 14800 -3730 14834 -3436
rect 14862 -3442 14920 -3436
rect 14862 -3706 14920 -3700
rect 15050 -3442 15108 -3436
rect 15050 -3706 15108 -3700
rect 15136 -3730 15170 -3436
rect 15198 -3442 15256 -3436
rect 15198 -3706 15256 -3700
rect 15386 -3442 15444 -3436
rect 15386 -3706 15444 -3700
rect 15472 -3730 15506 -3436
rect 15534 -3442 15592 -3436
rect 15534 -3706 15592 -3700
rect 15722 -3442 15780 -3436
rect 15722 -3706 15780 -3700
rect 15808 -3730 15842 -3436
rect 15870 -3442 15928 -3436
rect 15870 -3706 15928 -3700
rect 16058 -3442 16116 -3436
rect 16058 -3706 16116 -3700
rect 16144 -3730 16200 -3436
rect 14106 -4424 14128 -3736
rect 14162 -4424 14168 -3736
rect 14458 -3736 14504 -3730
rect 14106 -4558 14168 -4424
rect 14284 -4050 14342 -4040
rect 14284 -4436 14342 -4422
rect 14458 -4424 14464 -3736
rect 14498 -4424 14504 -3736
rect 14794 -3736 14840 -3730
rect 14458 -4558 14504 -4424
rect 14620 -4050 14678 -4040
rect 14620 -4436 14678 -4422
rect 14794 -4424 14800 -3736
rect 14834 -4424 14840 -3736
rect 15130 -3736 15176 -3730
rect 14794 -4558 14840 -4424
rect 14956 -4050 15014 -4040
rect 14956 -4436 15014 -4422
rect 15130 -4424 15136 -3736
rect 15170 -4424 15176 -3736
rect 15466 -3736 15512 -3730
rect 15130 -4558 15176 -4424
rect 15292 -4050 15350 -4040
rect 15292 -4436 15350 -4422
rect 15466 -4424 15472 -3736
rect 15506 -4424 15512 -3736
rect 15802 -3736 15848 -3730
rect 15466 -4558 15512 -4424
rect 15628 -4050 15686 -4040
rect 15628 -4436 15686 -4422
rect 15802 -4424 15808 -3736
rect 15842 -4424 15848 -3736
rect 16138 -3736 16200 -3730
rect 15802 -4558 15848 -4424
rect 15964 -4050 16022 -4040
rect 15964 -4436 16022 -4422
rect 16138 -4424 16144 -3736
rect 16178 -4424 16200 -3736
rect 16138 -4558 16200 -4424
rect 8712 -4616 8740 -4564
rect 9188 -4616 9216 -4564
rect 8712 -4646 9216 -4616
rect 14090 -4564 16214 -4558
rect 14090 -4616 14110 -4564
rect 16194 -4616 16214 -4564
rect 14090 -4622 16214 -4616
rect 16294 -4708 16406 -3160
rect 16294 -4876 16322 -4708
rect 16378 -4876 16406 -4708
rect 16294 -4886 16406 -4876
<< via1 >>
rect 13794 -1666 13850 -1498
rect 13924 -1820 16380 -1768
rect 14114 -2948 14172 -1972
rect 14518 -2948 14576 -1972
rect 14922 -2948 14980 -1972
rect 15326 -2948 15384 -1972
rect 15730 -2948 15788 -1972
rect 16134 -2948 16192 -1972
rect 14118 -3160 14342 -3108
rect 13764 -3300 13876 -3248
rect 14854 -3160 15078 -3108
rect 14480 -3300 14704 -3248
rect 15608 -3160 15832 -3108
rect 15234 -3300 15458 -3248
rect 15954 -3300 16178 -3248
rect 16294 -3160 16406 -3108
rect 9086 -4046 9198 -3756
rect 14190 -3700 14248 -3442
rect 14378 -3700 14436 -3442
rect 14526 -3700 14584 -3442
rect 14714 -3700 14772 -3442
rect 14862 -3700 14920 -3442
rect 15050 -3700 15108 -3442
rect 15198 -3700 15256 -3442
rect 15386 -3700 15444 -3442
rect 15534 -3700 15592 -3442
rect 15722 -3700 15780 -3442
rect 15870 -3700 15928 -3442
rect 16058 -3700 16116 -3442
rect 14284 -4422 14342 -4050
rect 14620 -4422 14678 -4050
rect 14956 -4422 15014 -4050
rect 15292 -4422 15350 -4050
rect 15628 -4422 15686 -4050
rect 15964 -4422 16022 -4050
rect 8740 -4616 9188 -4564
rect 14110 -4616 16194 -4564
rect 16322 -4876 16378 -4708
<< metal2 >>
rect 13764 -1498 13876 -1488
rect 13764 -1666 13794 -1498
rect 13850 -1666 13876 -1498
rect 13764 -1676 13876 -1666
rect 13904 -1768 20748 -1710
rect 13904 -1820 13924 -1768
rect 16380 -1820 20748 -1768
rect 13904 -1878 20748 -1820
rect 14114 -1972 14172 -1962
rect 14114 -2960 14172 -2948
rect 14518 -1972 14576 -1962
rect 14518 -2960 14576 -2948
rect 14922 -1972 14980 -1962
rect 14922 -2960 14980 -2948
rect 15326 -1972 15384 -1962
rect 15326 -2960 15384 -2948
rect 15730 -1972 15788 -1962
rect 15730 -2960 15788 -2948
rect 16134 -1972 16192 -1962
rect 16134 -2960 16192 -2948
rect 20524 -2250 20748 -1878
rect 14118 -3078 14240 -3050
rect 14040 -3108 16406 -3078
rect 14040 -3160 14118 -3108
rect 14342 -3160 14854 -3108
rect 15078 -3160 15608 -3108
rect 15832 -3160 16294 -3108
rect 14040 -3190 16406 -3160
rect 13764 -3248 16266 -3218
rect 13876 -3300 14480 -3248
rect 14704 -3300 15234 -3248
rect 15458 -3300 15954 -3248
rect 16178 -3300 16266 -3248
rect 13764 -3330 16266 -3300
rect 8712 -3442 16116 -3436
rect 8712 -3486 14190 -3442
rect 8712 -3598 8756 -3486
rect 9750 -3598 14190 -3486
rect 8712 -3660 14190 -3598
rect 14248 -3660 14378 -3442
rect 14190 -3706 14248 -3700
rect 14436 -3660 14526 -3442
rect 14378 -3706 14436 -3700
rect 14584 -3660 14714 -3442
rect 14526 -3706 14584 -3700
rect 14772 -3660 14862 -3442
rect 14714 -3706 14772 -3700
rect 14920 -3660 15050 -3442
rect 14862 -3706 14920 -3700
rect 15108 -3660 15198 -3442
rect 15050 -3706 15108 -3700
rect 15256 -3660 15386 -3442
rect 15198 -3706 15256 -3700
rect 15444 -3660 15534 -3442
rect 15386 -3706 15444 -3700
rect 15592 -3660 15722 -3442
rect 15534 -3706 15592 -3700
rect 15780 -3660 15870 -3442
rect 15722 -3706 15780 -3700
rect 15928 -3660 16058 -3442
rect 15870 -3706 15928 -3700
rect 16058 -3706 16116 -3700
rect 9078 -3756 9206 -3742
rect 9078 -4046 9086 -3756
rect 9198 -4046 9206 -3756
rect 9078 -4060 9206 -4046
rect 14284 -4050 14342 -4040
rect 14284 -4436 14342 -4422
rect 14620 -4050 14678 -4040
rect 14620 -4436 14678 -4422
rect 14956 -4050 15014 -4040
rect 14956 -4436 15014 -4422
rect 15292 -4050 15350 -4040
rect 15292 -4436 15350 -4422
rect 15628 -4050 15686 -4040
rect 15628 -4436 15686 -4422
rect 15964 -4050 16022 -4040
rect 20524 -4218 20580 -2250
rect 20692 -4218 20748 -2250
rect 20524 -4234 20748 -4218
rect 15964 -4436 16022 -4422
rect 8712 -4564 16214 -4534
rect 8712 -4616 8740 -4564
rect 9188 -4616 14110 -4564
rect 16194 -4616 16214 -4564
rect 8712 -4646 16214 -4616
rect 16294 -4708 16406 -4698
rect 16294 -4876 16322 -4708
rect 16378 -4876 16406 -4708
rect 16294 -4886 16406 -4876
<< via2 >>
rect 13794 -1666 13850 -1498
rect 14114 -2948 14172 -1972
rect 14518 -2948 14576 -1972
rect 14922 -2948 14980 -1972
rect 15326 -2948 15384 -1972
rect 15730 -2948 15788 -1972
rect 16134 -2948 16192 -1972
rect 8756 -3598 9750 -3486
rect 9086 -4046 9198 -3756
rect 14284 -4422 14342 -4050
rect 14620 -4422 14678 -4050
rect 14956 -4422 15014 -4050
rect 15292 -4422 15350 -4050
rect 15628 -4422 15686 -4050
rect 15964 -4422 16022 -4050
rect 20580 -4218 20692 -2250
rect 16322 -4876 16378 -4708
<< metal3 >>
rect 21292 5110 21532 5120
rect 21292 -790 21356 5110
rect 21468 -790 21532 5110
rect 8812 -1464 14892 -1454
rect 8812 -1498 15794 -1464
rect 8812 -1666 13794 -1498
rect 13850 -1666 15794 -1498
rect 8812 -1694 15794 -1666
rect 8712 -3486 9792 -1774
rect 8712 -3598 8756 -3486
rect 9750 -3598 9792 -3486
rect 8712 -3660 9792 -3598
rect 14108 -1972 14288 -1694
rect 14108 -2948 14114 -1972
rect 14172 -2948 14288 -1972
rect 14108 -3440 14288 -2948
rect 14512 -1972 14692 -1960
rect 14512 -2948 14518 -1972
rect 14576 -2948 14692 -1972
rect 9078 -3756 9206 -3742
rect 9078 -4046 9086 -3756
rect 9198 -4046 9206 -3756
rect 9078 -4060 9206 -4046
rect 14108 -4050 14348 -3440
rect 14108 -4422 14284 -4050
rect 14342 -4422 14348 -4050
rect 14108 -4428 14348 -4422
rect 14512 -4050 14692 -2948
rect 14512 -4422 14620 -4050
rect 14678 -4422 14692 -4050
rect 14512 -4682 14692 -4422
rect 14916 -1972 15096 -1694
rect 14916 -2948 14922 -1972
rect 14980 -2948 15096 -1972
rect 14916 -4050 15096 -2948
rect 14916 -4422 14956 -4050
rect 15014 -4422 15096 -4050
rect 14916 -4428 15096 -4422
rect 15270 -1972 15450 -1960
rect 15270 -2948 15326 -1972
rect 15384 -2948 15450 -1972
rect 15270 -4050 15450 -2948
rect 15270 -4422 15292 -4050
rect 15350 -4422 15450 -4050
rect 15270 -4682 15450 -4422
rect 15614 -1972 15794 -1694
rect 15614 -2948 15730 -1972
rect 15788 -2948 15794 -1972
rect 15614 -4050 15794 -2948
rect 15614 -4422 15628 -4050
rect 15686 -4422 15794 -4050
rect 15614 -4428 15794 -4422
rect 15958 -1972 16198 -1960
rect 15958 -2948 16134 -1972
rect 16192 -2948 16198 -1972
rect 21292 -2234 21532 -790
rect 15958 -2960 16198 -2948
rect 20524 -2250 21604 -2234
rect 15958 -4050 16144 -2960
rect 15958 -4422 15964 -4050
rect 16022 -4422 16144 -4050
rect 20524 -4218 20580 -2250
rect 20692 -4218 21604 -2250
rect 20524 -4234 21604 -4218
rect 15958 -4682 16144 -4422
rect 8812 -4708 16422 -4682
rect 8812 -4766 16322 -4708
rect 16378 -4766 16422 -4708
rect 8812 -4836 8818 -4766
rect 16416 -4836 16422 -4766
rect 8812 -4876 16322 -4836
rect 16378 -4876 16422 -4836
rect 8812 -4922 16422 -4876
rect 21292 -5384 21532 -4234
rect 21292 -11284 21356 -5384
rect 21468 -11284 21532 -5384
rect 21292 -11374 21532 -11284
<< via3 >>
rect 21356 -790 21468 5110
rect 9086 -4046 9198 -3756
rect 8818 -4836 16322 -4766
rect 16322 -4836 16378 -4766
rect 16378 -4836 16416 -4766
rect 21356 -11284 21468 -5384
<< metal4 >>
rect 8892 4816 14812 6008
rect 21132 5110 21474 5120
rect 21132 -790 21356 5110
rect 21468 -790 21474 5110
rect 21132 -800 21474 -790
rect 17956 -3706 18316 -1072
rect 9074 -3756 18316 -3706
rect 9074 -4046 9086 -3756
rect 9198 -4046 18316 -3756
rect 9074 -4066 18316 -4046
rect 8812 -4766 16422 -4760
rect 8812 -4836 8818 -4766
rect 16416 -4836 16422 -4766
rect 8812 -4942 16422 -4836
rect 8812 -5086 14892 -4942
rect 17956 -5092 18316 -4066
rect 21132 -5384 21474 -5374
rect 8892 -12474 14812 -11280
rect 21132 -11284 21356 -5384
rect 21468 -11284 21474 -5384
rect 21132 -11294 21474 -11284
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M11
timestamp 1681062556
transform 1 0 14266 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M12
timestamp 1681062556
transform 1 0 14360 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M13
timestamp 1681062556
transform 1 0 14938 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M14
timestamp 1681062556
transform 1 0 15032 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M15
timestamp 1681062556
transform 1 0 15610 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M16
timestamp 1681062556
transform 1 0 15704 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M21
timestamp 1681062556
transform 1 0 14602 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M22
timestamp 1681062556
transform 1 0 14696 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M23
timestamp 1681062556
transform 1 0 15274 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M24
timestamp 1681062556
transform 1 0 15368 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M25
timestamp 1681062556
transform 1 0 15946 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M26
timestamp 1681062556
transform 1 0 16040 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M31
timestamp 1681050310
transform 1 0 14079 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M32
timestamp 1681050310
transform 1 0 14207 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M33
timestamp 1681050310
transform 1 0 14887 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M34
timestamp 1681050310
transform 1 0 15015 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M35
timestamp 1681050310
transform 1 0 15695 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M36
timestamp 1681050310
transform 1 0 15823 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M41
timestamp 1681050310
transform 1 0 14483 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M42
timestamp 1681050310
transform 1 0 14611 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M43
timestamp 1681050310
transform 1 0 15291 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M44
timestamp 1681050310
transform 1 0 15419 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M45
timestamp 1681050310
transform 1 0 16099 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M46
timestamp 1681050310
transform 1 0 16227 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1680390383
transform 0 1 11852 -1 0 1722
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 1680390383
transform 0 1 11852 -1 0 -8188
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC31
timestamp 1680390383
transform 0 1 18172 -1 0 2014
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC32
timestamp 1680390383
transform 0 -1 18172 1 0 -8188
box -3186 -3040 3186 3040
<< labels >>
flabel metal3 8712 -3660 9792 -1774 0 FreeMono 1920 0 0 0 out1
port 2 nsew
flabel metal1 8712 -4646 9216 -3706 0 FreeMono 1280 0 0 0 vss
port 4 nsew
flabel metal3 20524 -4234 21604 -2234 0 FreeMono 1920 0 0 0 out2
port 3 nsew
flabel metal4 8892 -12474 14812 -11394 0 FreeMono 3200 0 0 0 vinn
port 1 nsew
flabel metal4 8892 4928 14812 6008 0 FreeMono 3200 0 0 0 vinp
port 0 nsew
<< end >>
