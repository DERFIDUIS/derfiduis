magic
tech sky130A
magscale 1 2
timestamp 1681683204
<< error_p >>
rect -29 141 29 147
rect -29 107 -17 141
rect -29 101 29 107
<< nmos >>
rect -18 -131 18 69
<< ndiff >>
rect -76 57 -18 69
rect -76 -119 -64 57
rect -30 -119 -18 57
rect -76 -131 -18 -119
rect 18 57 76 69
rect 18 -119 30 57
rect 64 -119 76 57
rect 18 -131 76 -119
<< ndiffc >>
rect -64 -119 -30 57
rect 30 -119 64 57
<< poly >>
rect -33 141 33 157
rect -33 107 -17 141
rect 17 107 33 141
rect -33 91 33 107
rect -18 69 18 91
rect -18 -157 18 -131
<< polycont >>
rect -17 107 17 141
<< locali >>
rect -33 107 -17 141
rect 17 107 33 141
rect -64 57 -30 73
rect -64 -135 -30 -119
rect 30 57 64 73
rect 30 -135 64 -119
<< viali >>
rect -17 107 17 141
rect -64 -119 -30 57
rect 30 -119 64 57
<< metal1 >>
rect -29 141 29 147
rect -29 107 -17 141
rect 17 107 29 141
rect -29 101 29 107
rect -70 57 -24 69
rect -70 -119 -64 57
rect -30 -119 -24 57
rect -70 -131 -24 -119
rect 24 57 70 69
rect 24 -119 30 57
rect 64 -119 70 57
rect 24 -131 70 -119
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
