** sch_path: /home/karlajcm/Documentos/TESIS DE
*+ GRADO/WORK_IN_PROGRESS/My_xschem/rectifier_lvt_01v8_tb.sch
**.subckt rectifier_lvt_01v8_tb vrec vinp vinn
*.iopin vrec
*.iopin vinp
*.iopin vinn
V1 vinp vinn sin(0 1 915000000 0 0)
.save i(v1)
x1 vinp vinn vrec GND rectifier
**** begin user architecture code

.control
save all
tran 0.5n 60u
plot vinp-vinn
plot vrec
.endc


** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

.include rectifier.spice

.GLOBAL GND
.end
