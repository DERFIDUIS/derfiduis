* NGSPICE file created from rectifier_lvt_01v8_initial.ext - technology: sky130A

.subckt rectifier_lvt_01v8_initial vinp vinn vss out2
M31 out2 vinn vinp out2 sky130_fd_pr__pfet_01v8_lvt ad=1.8e+13p pd=1.272e+08u as=4.35e+12p ps=3.174e+07u w=5e+06u l=350000u
M41 out2 vinp vinn out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=350000u
M11 vss vinn vinp vss sky130_fd_pr__nfet_01v8_lvt ad=1.8e+13p pd=1.272e+08u as=4.35e+12p ps=3.174e+07u w=5e+06u l=180000u
M12 vss vinn vinp vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M21 vss vinp vinn vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=4.35e+12p ps=3.174e+07u w=5e+06u l=180000u
M13 vinp vinn vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M42 out2 vinp vinn out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M22 vinn vinp vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M32 out2 vinn vinp out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M43 vinn vinp out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M14 vinp vinn vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M44 vinn vinp out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M23 vss vinp vinn vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M33 vinp vinn out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M24 vss vinp vinn vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M15 vss vinn vinp vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M16 vinp vinn vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M45 out2 vinp vinn out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M25 vinn vinp vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M34 out2 vinn vinp out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M26 vinn vinp vss vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=180000u
M46 vinn vinp out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M35 vinp vinn out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
M36 vinp vinn out2 out2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=350000u
.ends

