magic
tech sky130A
magscale 1 2
timestamp 1680252239
<< pwell >>
rect -201 -948 201 948
<< psubdiff >>
rect -165 878 -69 912
rect 69 878 165 912
rect -165 816 -131 878
rect 131 816 165 878
rect -165 -878 -131 -816
rect 131 -878 165 -816
rect -165 -912 -69 -878
rect 69 -912 165 -878
<< psubdiffcont >>
rect -69 878 69 912
rect -165 -816 -131 816
rect 131 -816 165 816
rect -69 -912 69 -878
<< xpolycontact >>
rect -35 350 35 782
rect -35 -782 35 -350
<< xpolyres >>
rect -35 -350 35 350
<< locali >>
rect -165 878 -69 912
rect 69 878 165 912
rect -165 816 -131 878
rect 131 816 165 878
rect -165 -878 -131 -816
rect 131 -878 165 -816
rect -165 -912 -69 -878
rect 69 -912 165 -878
<< viali >>
rect -19 367 19 764
rect -19 -764 19 -367
<< metal1 >>
rect -25 764 25 776
rect -25 367 -19 764
rect 19 367 25 764
rect -25 355 25 367
rect -25 -367 25 -355
rect -25 -764 -19 -367
rect 19 -764 25 -367
rect -25 -776 25 -764
<< res0p35 >>
rect -37 -352 37 352
<< properties >>
string FIXED_BBOX -148 -895 148 895
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 3.5 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 21.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
