** sch_path: /home/karlajcm/Documentos/TESIS DE
*+ GRADO/WORK_IN_PROGRESS/My_xschem/voltage_limiter_tb.sch
**.subckt voltage_limiter_tb vdd vrec
*.iopin vdd
*.iopin vrec
V1 vrec GND 1.8
.save i(v1)
x1 vrec vdd GND voltage_limiter
**** begin user architecture code

.control
save all
dc V1 0 6 0.1
plot vdd
.endc


** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  Documentos/TESIS DE GRADO/WORK_IN_PROGRESS/My_xschem/voltage_limiter.sym # of
*+ pins=3
** sym_path: /home/karlajcm/Documentos/TESIS DE GRADO/WORK_IN_PROGRESS/My_xschem/voltage_limiter.sym
** sch_path: /home/karlajcm/Documentos/TESIS DE GRADO/WORK_IN_PROGRESS/My_xschem/voltage_limiter.sch
.subckt voltage_limiter vrec vdd vss
*.iopin vss
*.iopin vrec
*.iopin vdd
XM4 net1 net4 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.7 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 vss net1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=16 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM2 net3 net3 net2 vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM3 net4 net4 net3 vdd sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XR3 vdd vrec vss sky130_fd_pr__res_xhigh_po W=1 L=2 mult=1 m=1
XR2 net1 vdd vss sky130_fd_pr__res_xhigh_po W=1 L=60 mult=1 m=1
XR4 vss net4 vss sky130_fd_pr__res_xhigh_po W=1 L=40 mult=1 m=1
.ends

.GLOBAL GND
.end
