** sch_path: /home/karlajcm/Documentos/TESIS DE
*+ GRADO/WORK_IN_PROGRESS/My_xschem/For_Layout/ring_oscillator.sch
.subckt ring_oscillator vtemp vss vdd vosc
*.PININFO vtemp:B vss:B vdd:B vosc:B
M1 net1 vosc vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=12 nf=1 m=1
M2 net1 vosc vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=4 nf=1 m=1
M3 net2 net1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=12 nf=1 m=1
M4 net2 net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=4 nf=1 m=1
M5 vosc net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=12 nf=1 m=1
M6 vosc net2 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=4 nf=1 m=1
XC1 vosc vtemp vss sky130_fd_pr__cap_var_lvt W=5 L=5 VM=1 m=1
XC2 net2 vtemp vss sky130_fd_pr__cap_var_lvt W=5 L=5 VM=1 m=1
XC3 net1 vtemp vss sky130_fd_pr__cap_var_lvt W=5 L=5 VM=1 m=1
.ends
.end
