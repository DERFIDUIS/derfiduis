magic
tech sky130A
magscale 1 2
timestamp 1681253575
<< nwell >>
rect 10966 -3060 11032 -1898
rect 11370 -3060 11484 -1898
rect 11774 -3060 11888 -1898
rect 12178 -3060 12292 -1898
rect 12582 -3060 12696 -1898
rect 12986 -3060 13100 -1898
rect 13438 -3060 13504 -1898
<< ndiff >>
rect 11270 -4436 11272 -3436
rect 11518 -4436 11520 -3436
rect 11606 -4436 11608 -3436
rect 11854 -4436 11856 -3436
rect 11942 -4436 11944 -3436
rect 12190 -4436 12192 -3436
rect 12278 -4436 12280 -3436
rect 12526 -4436 12528 -3436
rect 12614 -4436 12616 -3436
rect 12862 -4436 12864 -3436
rect 12950 -4436 12952 -3436
rect 13198 -4436 13200 -3436
<< pdiff >>
rect 11066 -2960 11068 -1960
rect 11382 -2960 11384 -1960
rect 11470 -2960 11472 -1960
rect 11786 -2960 11788 -1960
rect 11874 -2960 11876 -1960
rect 12190 -2960 12192 -1960
rect 12278 -2960 12280 -1960
rect 12594 -2960 12596 -1960
rect 12682 -2960 12684 -1960
rect 12998 -2960 13000 -1960
rect 13086 -2960 13088 -1960
rect 13402 -2960 13404 -1960
<< psubdiff >>
rect 11206 -3490 11270 -3436
rect 11206 -3524 11210 -3490
rect 11244 -3524 11270 -3490
rect 11206 -3558 11270 -3524
rect 11206 -3592 11210 -3558
rect 11244 -3592 11270 -3558
rect 11206 -3626 11270 -3592
rect 11206 -3660 11210 -3626
rect 11244 -3660 11270 -3626
rect 11206 -3694 11270 -3660
rect 11206 -3728 11210 -3694
rect 11244 -3728 11270 -3694
rect 11206 -3762 11270 -3728
rect 11206 -3796 11210 -3762
rect 11244 -3796 11270 -3762
rect 11206 -3830 11270 -3796
rect 11206 -3864 11210 -3830
rect 11244 -3864 11270 -3830
rect 11206 -3898 11270 -3864
rect 11206 -3932 11210 -3898
rect 11244 -3932 11270 -3898
rect 11206 -3966 11270 -3932
rect 11206 -4000 11210 -3966
rect 11244 -4000 11270 -3966
rect 11206 -4034 11270 -4000
rect 11206 -4068 11210 -4034
rect 11244 -4068 11270 -4034
rect 11206 -4102 11270 -4068
rect 11206 -4136 11210 -4102
rect 11244 -4136 11270 -4102
rect 11206 -4170 11270 -4136
rect 11206 -4204 11210 -4170
rect 11244 -4204 11270 -4170
rect 11206 -4238 11270 -4204
rect 11206 -4272 11210 -4238
rect 11244 -4272 11270 -4238
rect 11206 -4306 11270 -4272
rect 11206 -4340 11210 -4306
rect 11244 -4340 11270 -4306
rect 11206 -4374 11270 -4340
rect 11206 -4408 11210 -4374
rect 11244 -4408 11270 -4374
rect 11206 -4436 11270 -4408
rect 11520 -3464 11606 -3436
rect 11520 -3498 11546 -3464
rect 11580 -3498 11606 -3464
rect 11520 -3532 11606 -3498
rect 11520 -3566 11546 -3532
rect 11580 -3566 11606 -3532
rect 11520 -3600 11606 -3566
rect 11520 -3634 11546 -3600
rect 11580 -3634 11606 -3600
rect 11520 -3668 11606 -3634
rect 11520 -3702 11546 -3668
rect 11580 -3702 11606 -3668
rect 11520 -3736 11606 -3702
rect 11520 -3770 11546 -3736
rect 11580 -3770 11606 -3736
rect 11520 -3804 11606 -3770
rect 11520 -3838 11546 -3804
rect 11580 -3838 11606 -3804
rect 11520 -3872 11606 -3838
rect 11520 -3906 11546 -3872
rect 11580 -3906 11606 -3872
rect 11520 -3940 11606 -3906
rect 11520 -3974 11546 -3940
rect 11580 -3974 11606 -3940
rect 11520 -4008 11606 -3974
rect 11520 -4042 11546 -4008
rect 11580 -4042 11606 -4008
rect 11520 -4076 11606 -4042
rect 11520 -4110 11546 -4076
rect 11580 -4110 11606 -4076
rect 11520 -4144 11606 -4110
rect 11520 -4178 11546 -4144
rect 11580 -4178 11606 -4144
rect 11520 -4212 11606 -4178
rect 11520 -4246 11546 -4212
rect 11580 -4246 11606 -4212
rect 11520 -4280 11606 -4246
rect 11520 -4314 11546 -4280
rect 11580 -4314 11606 -4280
rect 11520 -4348 11606 -4314
rect 11520 -4382 11546 -4348
rect 11580 -4382 11606 -4348
rect 11520 -4436 11606 -4382
rect 11856 -3464 11942 -3436
rect 11856 -3498 11882 -3464
rect 11916 -3498 11942 -3464
rect 11856 -3532 11942 -3498
rect 11856 -3566 11882 -3532
rect 11916 -3566 11942 -3532
rect 11856 -3600 11942 -3566
rect 11856 -3634 11882 -3600
rect 11916 -3634 11942 -3600
rect 11856 -3668 11942 -3634
rect 11856 -3702 11882 -3668
rect 11916 -3702 11942 -3668
rect 11856 -3736 11942 -3702
rect 11856 -3770 11882 -3736
rect 11916 -3770 11942 -3736
rect 11856 -3804 11942 -3770
rect 11856 -3838 11882 -3804
rect 11916 -3838 11942 -3804
rect 11856 -3872 11942 -3838
rect 11856 -3906 11882 -3872
rect 11916 -3906 11942 -3872
rect 11856 -3940 11942 -3906
rect 11856 -3974 11882 -3940
rect 11916 -3974 11942 -3940
rect 11856 -4008 11942 -3974
rect 11856 -4042 11882 -4008
rect 11916 -4042 11942 -4008
rect 11856 -4076 11942 -4042
rect 11856 -4110 11882 -4076
rect 11916 -4110 11942 -4076
rect 11856 -4144 11942 -4110
rect 11856 -4178 11882 -4144
rect 11916 -4178 11942 -4144
rect 11856 -4212 11942 -4178
rect 11856 -4246 11882 -4212
rect 11916 -4246 11942 -4212
rect 11856 -4280 11942 -4246
rect 11856 -4314 11882 -4280
rect 11916 -4314 11942 -4280
rect 11856 -4348 11942 -4314
rect 11856 -4382 11882 -4348
rect 11916 -4382 11942 -4348
rect 11856 -4436 11942 -4382
rect 12192 -3464 12278 -3436
rect 12192 -3498 12218 -3464
rect 12252 -3498 12278 -3464
rect 12192 -3532 12278 -3498
rect 12192 -3566 12218 -3532
rect 12252 -3566 12278 -3532
rect 12192 -3600 12278 -3566
rect 12192 -3634 12218 -3600
rect 12252 -3634 12278 -3600
rect 12192 -3668 12278 -3634
rect 12192 -3702 12218 -3668
rect 12252 -3702 12278 -3668
rect 12192 -3736 12278 -3702
rect 12192 -3770 12218 -3736
rect 12252 -3770 12278 -3736
rect 12192 -3804 12278 -3770
rect 12192 -3838 12218 -3804
rect 12252 -3838 12278 -3804
rect 12192 -3872 12278 -3838
rect 12192 -3906 12218 -3872
rect 12252 -3906 12278 -3872
rect 12192 -3940 12278 -3906
rect 12192 -3974 12218 -3940
rect 12252 -3974 12278 -3940
rect 12192 -4008 12278 -3974
rect 12192 -4042 12218 -4008
rect 12252 -4042 12278 -4008
rect 12192 -4076 12278 -4042
rect 12192 -4110 12218 -4076
rect 12252 -4110 12278 -4076
rect 12192 -4144 12278 -4110
rect 12192 -4178 12218 -4144
rect 12252 -4178 12278 -4144
rect 12192 -4212 12278 -4178
rect 12192 -4246 12218 -4212
rect 12252 -4246 12278 -4212
rect 12192 -4280 12278 -4246
rect 12192 -4314 12218 -4280
rect 12252 -4314 12278 -4280
rect 12192 -4348 12278 -4314
rect 12192 -4382 12218 -4348
rect 12252 -4382 12278 -4348
rect 12192 -4436 12278 -4382
rect 12528 -3464 12614 -3436
rect 12528 -3498 12554 -3464
rect 12588 -3498 12614 -3464
rect 12528 -3532 12614 -3498
rect 12528 -3566 12554 -3532
rect 12588 -3566 12614 -3532
rect 12528 -3600 12614 -3566
rect 12528 -3634 12554 -3600
rect 12588 -3634 12614 -3600
rect 12528 -3668 12614 -3634
rect 12528 -3702 12554 -3668
rect 12588 -3702 12614 -3668
rect 12528 -3736 12614 -3702
rect 12528 -3770 12554 -3736
rect 12588 -3770 12614 -3736
rect 12528 -3804 12614 -3770
rect 12528 -3838 12554 -3804
rect 12588 -3838 12614 -3804
rect 12528 -3872 12614 -3838
rect 12528 -3906 12554 -3872
rect 12588 -3906 12614 -3872
rect 12528 -3940 12614 -3906
rect 12528 -3974 12554 -3940
rect 12588 -3974 12614 -3940
rect 12528 -4008 12614 -3974
rect 12528 -4042 12554 -4008
rect 12588 -4042 12614 -4008
rect 12528 -4076 12614 -4042
rect 12528 -4110 12554 -4076
rect 12588 -4110 12614 -4076
rect 12528 -4144 12614 -4110
rect 12528 -4178 12554 -4144
rect 12588 -4178 12614 -4144
rect 12528 -4212 12614 -4178
rect 12528 -4246 12554 -4212
rect 12588 -4246 12614 -4212
rect 12528 -4280 12614 -4246
rect 12528 -4314 12554 -4280
rect 12588 -4314 12614 -4280
rect 12528 -4348 12614 -4314
rect 12528 -4382 12554 -4348
rect 12588 -4382 12614 -4348
rect 12528 -4436 12614 -4382
rect 12864 -3464 12950 -3436
rect 12864 -3498 12890 -3464
rect 12924 -3498 12950 -3464
rect 12864 -3532 12950 -3498
rect 12864 -3566 12890 -3532
rect 12924 -3566 12950 -3532
rect 12864 -3600 12950 -3566
rect 12864 -3634 12890 -3600
rect 12924 -3634 12950 -3600
rect 12864 -3668 12950 -3634
rect 12864 -3702 12890 -3668
rect 12924 -3702 12950 -3668
rect 12864 -3736 12950 -3702
rect 12864 -3770 12890 -3736
rect 12924 -3770 12950 -3736
rect 12864 -3804 12950 -3770
rect 12864 -3838 12890 -3804
rect 12924 -3838 12950 -3804
rect 12864 -3872 12950 -3838
rect 12864 -3906 12890 -3872
rect 12924 -3906 12950 -3872
rect 12864 -3940 12950 -3906
rect 12864 -3974 12890 -3940
rect 12924 -3974 12950 -3940
rect 12864 -4008 12950 -3974
rect 12864 -4042 12890 -4008
rect 12924 -4042 12950 -4008
rect 12864 -4076 12950 -4042
rect 12864 -4110 12890 -4076
rect 12924 -4110 12950 -4076
rect 12864 -4144 12950 -4110
rect 12864 -4178 12890 -4144
rect 12924 -4178 12950 -4144
rect 12864 -4212 12950 -4178
rect 12864 -4246 12890 -4212
rect 12924 -4246 12950 -4212
rect 12864 -4280 12950 -4246
rect 12864 -4314 12890 -4280
rect 12924 -4314 12950 -4280
rect 12864 -4348 12950 -4314
rect 12864 -4382 12890 -4348
rect 12924 -4382 12950 -4348
rect 12864 -4436 12950 -4382
rect 13200 -3464 13264 -3436
rect 13200 -3498 13226 -3464
rect 13260 -3498 13264 -3464
rect 13200 -3532 13264 -3498
rect 13200 -3566 13226 -3532
rect 13260 -3566 13264 -3532
rect 13200 -3600 13264 -3566
rect 13200 -3634 13226 -3600
rect 13260 -3634 13264 -3600
rect 13200 -3668 13264 -3634
rect 13200 -3702 13226 -3668
rect 13260 -3702 13264 -3668
rect 13200 -3736 13264 -3702
rect 13200 -3770 13226 -3736
rect 13260 -3770 13264 -3736
rect 13200 -3804 13264 -3770
rect 13200 -3838 13226 -3804
rect 13260 -3838 13264 -3804
rect 13200 -3872 13264 -3838
rect 13200 -3906 13226 -3872
rect 13260 -3906 13264 -3872
rect 13200 -3940 13264 -3906
rect 13200 -3974 13226 -3940
rect 13260 -3974 13264 -3940
rect 13200 -4008 13264 -3974
rect 13200 -4042 13226 -4008
rect 13260 -4042 13264 -4008
rect 13200 -4076 13264 -4042
rect 13200 -4110 13226 -4076
rect 13260 -4110 13264 -4076
rect 13200 -4144 13264 -4110
rect 13200 -4178 13226 -4144
rect 13260 -4178 13264 -4144
rect 13200 -4212 13264 -4178
rect 13200 -4246 13226 -4212
rect 13260 -4246 13264 -4212
rect 13200 -4280 13264 -4246
rect 13200 -4314 13226 -4280
rect 13260 -4314 13264 -4280
rect 13200 -4348 13264 -4314
rect 13200 -4382 13226 -4348
rect 13260 -4382 13264 -4348
rect 13200 -4436 13264 -4382
<< nsubdiff >>
rect 11002 -2014 11066 -1960
rect 11002 -2048 11006 -2014
rect 11040 -2048 11066 -2014
rect 11002 -2082 11066 -2048
rect 11002 -2116 11006 -2082
rect 11040 -2116 11066 -2082
rect 11002 -2150 11066 -2116
rect 11002 -2184 11006 -2150
rect 11040 -2184 11066 -2150
rect 11002 -2218 11066 -2184
rect 11002 -2252 11006 -2218
rect 11040 -2252 11066 -2218
rect 11002 -2286 11066 -2252
rect 11002 -2320 11006 -2286
rect 11040 -2320 11066 -2286
rect 11002 -2354 11066 -2320
rect 11002 -2388 11006 -2354
rect 11040 -2388 11066 -2354
rect 11002 -2422 11066 -2388
rect 11002 -2456 11006 -2422
rect 11040 -2456 11066 -2422
rect 11002 -2490 11066 -2456
rect 11002 -2524 11006 -2490
rect 11040 -2524 11066 -2490
rect 11002 -2558 11066 -2524
rect 11002 -2592 11006 -2558
rect 11040 -2592 11066 -2558
rect 11002 -2626 11066 -2592
rect 11002 -2660 11006 -2626
rect 11040 -2660 11066 -2626
rect 11002 -2694 11066 -2660
rect 11002 -2728 11006 -2694
rect 11040 -2728 11066 -2694
rect 11002 -2762 11066 -2728
rect 11002 -2796 11006 -2762
rect 11040 -2796 11066 -2762
rect 11002 -2830 11066 -2796
rect 11002 -2864 11006 -2830
rect 11040 -2864 11066 -2830
rect 11002 -2898 11066 -2864
rect 11002 -2932 11006 -2898
rect 11040 -2932 11066 -2898
rect 11002 -2960 11066 -2932
rect 11384 -1988 11470 -1960
rect 11384 -2022 11410 -1988
rect 11444 -2022 11470 -1988
rect 11384 -2056 11470 -2022
rect 11384 -2090 11410 -2056
rect 11444 -2090 11470 -2056
rect 11384 -2124 11470 -2090
rect 11384 -2158 11410 -2124
rect 11444 -2158 11470 -2124
rect 11384 -2192 11470 -2158
rect 11384 -2226 11410 -2192
rect 11444 -2226 11470 -2192
rect 11384 -2260 11470 -2226
rect 11384 -2294 11410 -2260
rect 11444 -2294 11470 -2260
rect 11384 -2328 11470 -2294
rect 11384 -2362 11410 -2328
rect 11444 -2362 11470 -2328
rect 11384 -2396 11470 -2362
rect 11384 -2430 11410 -2396
rect 11444 -2430 11470 -2396
rect 11384 -2464 11470 -2430
rect 11384 -2498 11410 -2464
rect 11444 -2498 11470 -2464
rect 11384 -2532 11470 -2498
rect 11384 -2566 11410 -2532
rect 11444 -2566 11470 -2532
rect 11384 -2600 11470 -2566
rect 11384 -2634 11410 -2600
rect 11444 -2634 11470 -2600
rect 11384 -2668 11470 -2634
rect 11384 -2702 11410 -2668
rect 11444 -2702 11470 -2668
rect 11384 -2736 11470 -2702
rect 11384 -2770 11410 -2736
rect 11444 -2770 11470 -2736
rect 11384 -2804 11470 -2770
rect 11384 -2838 11410 -2804
rect 11444 -2838 11470 -2804
rect 11384 -2872 11470 -2838
rect 11384 -2906 11410 -2872
rect 11444 -2906 11470 -2872
rect 11384 -2960 11470 -2906
rect 11788 -1988 11874 -1960
rect 11788 -2022 11814 -1988
rect 11848 -2022 11874 -1988
rect 11788 -2056 11874 -2022
rect 11788 -2090 11814 -2056
rect 11848 -2090 11874 -2056
rect 11788 -2124 11874 -2090
rect 11788 -2158 11814 -2124
rect 11848 -2158 11874 -2124
rect 11788 -2192 11874 -2158
rect 11788 -2226 11814 -2192
rect 11848 -2226 11874 -2192
rect 11788 -2260 11874 -2226
rect 11788 -2294 11814 -2260
rect 11848 -2294 11874 -2260
rect 11788 -2328 11874 -2294
rect 11788 -2362 11814 -2328
rect 11848 -2362 11874 -2328
rect 11788 -2396 11874 -2362
rect 11788 -2430 11814 -2396
rect 11848 -2430 11874 -2396
rect 11788 -2464 11874 -2430
rect 11788 -2498 11814 -2464
rect 11848 -2498 11874 -2464
rect 11788 -2532 11874 -2498
rect 11788 -2566 11814 -2532
rect 11848 -2566 11874 -2532
rect 11788 -2600 11874 -2566
rect 11788 -2634 11814 -2600
rect 11848 -2634 11874 -2600
rect 11788 -2668 11874 -2634
rect 11788 -2702 11814 -2668
rect 11848 -2702 11874 -2668
rect 11788 -2736 11874 -2702
rect 11788 -2770 11814 -2736
rect 11848 -2770 11874 -2736
rect 11788 -2804 11874 -2770
rect 11788 -2838 11814 -2804
rect 11848 -2838 11874 -2804
rect 11788 -2872 11874 -2838
rect 11788 -2906 11814 -2872
rect 11848 -2906 11874 -2872
rect 11788 -2960 11874 -2906
rect 12192 -1988 12278 -1960
rect 12192 -2022 12218 -1988
rect 12252 -2022 12278 -1988
rect 12192 -2056 12278 -2022
rect 12192 -2090 12218 -2056
rect 12252 -2090 12278 -2056
rect 12192 -2124 12278 -2090
rect 12192 -2158 12218 -2124
rect 12252 -2158 12278 -2124
rect 12192 -2192 12278 -2158
rect 12192 -2226 12218 -2192
rect 12252 -2226 12278 -2192
rect 12192 -2260 12278 -2226
rect 12192 -2294 12218 -2260
rect 12252 -2294 12278 -2260
rect 12192 -2328 12278 -2294
rect 12192 -2362 12218 -2328
rect 12252 -2362 12278 -2328
rect 12192 -2396 12278 -2362
rect 12192 -2430 12218 -2396
rect 12252 -2430 12278 -2396
rect 12192 -2464 12278 -2430
rect 12192 -2498 12218 -2464
rect 12252 -2498 12278 -2464
rect 12192 -2532 12278 -2498
rect 12192 -2566 12218 -2532
rect 12252 -2566 12278 -2532
rect 12192 -2600 12278 -2566
rect 12192 -2634 12218 -2600
rect 12252 -2634 12278 -2600
rect 12192 -2668 12278 -2634
rect 12192 -2702 12218 -2668
rect 12252 -2702 12278 -2668
rect 12192 -2736 12278 -2702
rect 12192 -2770 12218 -2736
rect 12252 -2770 12278 -2736
rect 12192 -2804 12278 -2770
rect 12192 -2838 12218 -2804
rect 12252 -2838 12278 -2804
rect 12192 -2872 12278 -2838
rect 12192 -2906 12218 -2872
rect 12252 -2906 12278 -2872
rect 12192 -2960 12278 -2906
rect 12596 -1988 12682 -1960
rect 12596 -2022 12622 -1988
rect 12656 -2022 12682 -1988
rect 12596 -2056 12682 -2022
rect 12596 -2090 12622 -2056
rect 12656 -2090 12682 -2056
rect 12596 -2124 12682 -2090
rect 12596 -2158 12622 -2124
rect 12656 -2158 12682 -2124
rect 12596 -2192 12682 -2158
rect 12596 -2226 12622 -2192
rect 12656 -2226 12682 -2192
rect 12596 -2260 12682 -2226
rect 12596 -2294 12622 -2260
rect 12656 -2294 12682 -2260
rect 12596 -2328 12682 -2294
rect 12596 -2362 12622 -2328
rect 12656 -2362 12682 -2328
rect 12596 -2396 12682 -2362
rect 12596 -2430 12622 -2396
rect 12656 -2430 12682 -2396
rect 12596 -2464 12682 -2430
rect 12596 -2498 12622 -2464
rect 12656 -2498 12682 -2464
rect 12596 -2532 12682 -2498
rect 12596 -2566 12622 -2532
rect 12656 -2566 12682 -2532
rect 12596 -2600 12682 -2566
rect 12596 -2634 12622 -2600
rect 12656 -2634 12682 -2600
rect 12596 -2668 12682 -2634
rect 12596 -2702 12622 -2668
rect 12656 -2702 12682 -2668
rect 12596 -2736 12682 -2702
rect 12596 -2770 12622 -2736
rect 12656 -2770 12682 -2736
rect 12596 -2804 12682 -2770
rect 12596 -2838 12622 -2804
rect 12656 -2838 12682 -2804
rect 12596 -2872 12682 -2838
rect 12596 -2906 12622 -2872
rect 12656 -2906 12682 -2872
rect 12596 -2960 12682 -2906
rect 13000 -1988 13086 -1960
rect 13000 -2022 13026 -1988
rect 13060 -2022 13086 -1988
rect 13000 -2056 13086 -2022
rect 13000 -2090 13026 -2056
rect 13060 -2090 13086 -2056
rect 13000 -2124 13086 -2090
rect 13000 -2158 13026 -2124
rect 13060 -2158 13086 -2124
rect 13000 -2192 13086 -2158
rect 13000 -2226 13026 -2192
rect 13060 -2226 13086 -2192
rect 13000 -2260 13086 -2226
rect 13000 -2294 13026 -2260
rect 13060 -2294 13086 -2260
rect 13000 -2328 13086 -2294
rect 13000 -2362 13026 -2328
rect 13060 -2362 13086 -2328
rect 13000 -2396 13086 -2362
rect 13000 -2430 13026 -2396
rect 13060 -2430 13086 -2396
rect 13000 -2464 13086 -2430
rect 13000 -2498 13026 -2464
rect 13060 -2498 13086 -2464
rect 13000 -2532 13086 -2498
rect 13000 -2566 13026 -2532
rect 13060 -2566 13086 -2532
rect 13000 -2600 13086 -2566
rect 13000 -2634 13026 -2600
rect 13060 -2634 13086 -2600
rect 13000 -2668 13086 -2634
rect 13000 -2702 13026 -2668
rect 13060 -2702 13086 -2668
rect 13000 -2736 13086 -2702
rect 13000 -2770 13026 -2736
rect 13060 -2770 13086 -2736
rect 13000 -2804 13086 -2770
rect 13000 -2838 13026 -2804
rect 13060 -2838 13086 -2804
rect 13000 -2872 13086 -2838
rect 13000 -2906 13026 -2872
rect 13060 -2906 13086 -2872
rect 13000 -2960 13086 -2906
rect 13404 -1988 13468 -1960
rect 13404 -2022 13430 -1988
rect 13464 -2022 13468 -1988
rect 13404 -2056 13468 -2022
rect 13404 -2090 13430 -2056
rect 13464 -2090 13468 -2056
rect 13404 -2124 13468 -2090
rect 13404 -2158 13430 -2124
rect 13464 -2158 13468 -2124
rect 13404 -2192 13468 -2158
rect 13404 -2226 13430 -2192
rect 13464 -2226 13468 -2192
rect 13404 -2260 13468 -2226
rect 13404 -2294 13430 -2260
rect 13464 -2294 13468 -2260
rect 13404 -2328 13468 -2294
rect 13404 -2362 13430 -2328
rect 13464 -2362 13468 -2328
rect 13404 -2396 13468 -2362
rect 13404 -2430 13430 -2396
rect 13464 -2430 13468 -2396
rect 13404 -2464 13468 -2430
rect 13404 -2498 13430 -2464
rect 13464 -2498 13468 -2464
rect 13404 -2532 13468 -2498
rect 13404 -2566 13430 -2532
rect 13464 -2566 13468 -2532
rect 13404 -2600 13468 -2566
rect 13404 -2634 13430 -2600
rect 13464 -2634 13468 -2600
rect 13404 -2668 13468 -2634
rect 13404 -2702 13430 -2668
rect 13464 -2702 13468 -2668
rect 13404 -2736 13468 -2702
rect 13404 -2770 13430 -2736
rect 13464 -2770 13468 -2736
rect 13404 -2804 13468 -2770
rect 13404 -2838 13430 -2804
rect 13464 -2838 13468 -2804
rect 13404 -2872 13468 -2838
rect 13404 -2906 13430 -2872
rect 13464 -2906 13468 -2872
rect 13404 -2960 13468 -2906
<< psubdiffcont >>
rect 11210 -3524 11244 -3490
rect 11210 -3592 11244 -3558
rect 11210 -3660 11244 -3626
rect 11210 -3728 11244 -3694
rect 11210 -3796 11244 -3762
rect 11210 -3864 11244 -3830
rect 11210 -3932 11244 -3898
rect 11210 -4000 11244 -3966
rect 11210 -4068 11244 -4034
rect 11210 -4136 11244 -4102
rect 11210 -4204 11244 -4170
rect 11210 -4272 11244 -4238
rect 11210 -4340 11244 -4306
rect 11210 -4408 11244 -4374
rect 11546 -3498 11580 -3464
rect 11546 -3566 11580 -3532
rect 11546 -3634 11580 -3600
rect 11546 -3702 11580 -3668
rect 11546 -3770 11580 -3736
rect 11546 -3838 11580 -3804
rect 11546 -3906 11580 -3872
rect 11546 -3974 11580 -3940
rect 11546 -4042 11580 -4008
rect 11546 -4110 11580 -4076
rect 11546 -4178 11580 -4144
rect 11546 -4246 11580 -4212
rect 11546 -4314 11580 -4280
rect 11546 -4382 11580 -4348
rect 11882 -3498 11916 -3464
rect 11882 -3566 11916 -3532
rect 11882 -3634 11916 -3600
rect 11882 -3702 11916 -3668
rect 11882 -3770 11916 -3736
rect 11882 -3838 11916 -3804
rect 11882 -3906 11916 -3872
rect 11882 -3974 11916 -3940
rect 11882 -4042 11916 -4008
rect 11882 -4110 11916 -4076
rect 11882 -4178 11916 -4144
rect 11882 -4246 11916 -4212
rect 11882 -4314 11916 -4280
rect 11882 -4382 11916 -4348
rect 12218 -3498 12252 -3464
rect 12218 -3566 12252 -3532
rect 12218 -3634 12252 -3600
rect 12218 -3702 12252 -3668
rect 12218 -3770 12252 -3736
rect 12218 -3838 12252 -3804
rect 12218 -3906 12252 -3872
rect 12218 -3974 12252 -3940
rect 12218 -4042 12252 -4008
rect 12218 -4110 12252 -4076
rect 12218 -4178 12252 -4144
rect 12218 -4246 12252 -4212
rect 12218 -4314 12252 -4280
rect 12218 -4382 12252 -4348
rect 12554 -3498 12588 -3464
rect 12554 -3566 12588 -3532
rect 12554 -3634 12588 -3600
rect 12554 -3702 12588 -3668
rect 12554 -3770 12588 -3736
rect 12554 -3838 12588 -3804
rect 12554 -3906 12588 -3872
rect 12554 -3974 12588 -3940
rect 12554 -4042 12588 -4008
rect 12554 -4110 12588 -4076
rect 12554 -4178 12588 -4144
rect 12554 -4246 12588 -4212
rect 12554 -4314 12588 -4280
rect 12554 -4382 12588 -4348
rect 12890 -3498 12924 -3464
rect 12890 -3566 12924 -3532
rect 12890 -3634 12924 -3600
rect 12890 -3702 12924 -3668
rect 12890 -3770 12924 -3736
rect 12890 -3838 12924 -3804
rect 12890 -3906 12924 -3872
rect 12890 -3974 12924 -3940
rect 12890 -4042 12924 -4008
rect 12890 -4110 12924 -4076
rect 12890 -4178 12924 -4144
rect 12890 -4246 12924 -4212
rect 12890 -4314 12924 -4280
rect 12890 -4382 12924 -4348
rect 13226 -3498 13260 -3464
rect 13226 -3566 13260 -3532
rect 13226 -3634 13260 -3600
rect 13226 -3702 13260 -3668
rect 13226 -3770 13260 -3736
rect 13226 -3838 13260 -3804
rect 13226 -3906 13260 -3872
rect 13226 -3974 13260 -3940
rect 13226 -4042 13260 -4008
rect 13226 -4110 13260 -4076
rect 13226 -4178 13260 -4144
rect 13226 -4246 13260 -4212
rect 13226 -4314 13260 -4280
rect 13226 -4382 13260 -4348
<< nsubdiffcont >>
rect 11006 -2048 11040 -2014
rect 11006 -2116 11040 -2082
rect 11006 -2184 11040 -2150
rect 11006 -2252 11040 -2218
rect 11006 -2320 11040 -2286
rect 11006 -2388 11040 -2354
rect 11006 -2456 11040 -2422
rect 11006 -2524 11040 -2490
rect 11006 -2592 11040 -2558
rect 11006 -2660 11040 -2626
rect 11006 -2728 11040 -2694
rect 11006 -2796 11040 -2762
rect 11006 -2864 11040 -2830
rect 11006 -2932 11040 -2898
rect 11410 -2022 11444 -1988
rect 11410 -2090 11444 -2056
rect 11410 -2158 11444 -2124
rect 11410 -2226 11444 -2192
rect 11410 -2294 11444 -2260
rect 11410 -2362 11444 -2328
rect 11410 -2430 11444 -2396
rect 11410 -2498 11444 -2464
rect 11410 -2566 11444 -2532
rect 11410 -2634 11444 -2600
rect 11410 -2702 11444 -2668
rect 11410 -2770 11444 -2736
rect 11410 -2838 11444 -2804
rect 11410 -2906 11444 -2872
rect 11814 -2022 11848 -1988
rect 11814 -2090 11848 -2056
rect 11814 -2158 11848 -2124
rect 11814 -2226 11848 -2192
rect 11814 -2294 11848 -2260
rect 11814 -2362 11848 -2328
rect 11814 -2430 11848 -2396
rect 11814 -2498 11848 -2464
rect 11814 -2566 11848 -2532
rect 11814 -2634 11848 -2600
rect 11814 -2702 11848 -2668
rect 11814 -2770 11848 -2736
rect 11814 -2838 11848 -2804
rect 11814 -2906 11848 -2872
rect 12218 -2022 12252 -1988
rect 12218 -2090 12252 -2056
rect 12218 -2158 12252 -2124
rect 12218 -2226 12252 -2192
rect 12218 -2294 12252 -2260
rect 12218 -2362 12252 -2328
rect 12218 -2430 12252 -2396
rect 12218 -2498 12252 -2464
rect 12218 -2566 12252 -2532
rect 12218 -2634 12252 -2600
rect 12218 -2702 12252 -2668
rect 12218 -2770 12252 -2736
rect 12218 -2838 12252 -2804
rect 12218 -2906 12252 -2872
rect 12622 -2022 12656 -1988
rect 12622 -2090 12656 -2056
rect 12622 -2158 12656 -2124
rect 12622 -2226 12656 -2192
rect 12622 -2294 12656 -2260
rect 12622 -2362 12656 -2328
rect 12622 -2430 12656 -2396
rect 12622 -2498 12656 -2464
rect 12622 -2566 12656 -2532
rect 12622 -2634 12656 -2600
rect 12622 -2702 12656 -2668
rect 12622 -2770 12656 -2736
rect 12622 -2838 12656 -2804
rect 12622 -2906 12656 -2872
rect 13026 -2022 13060 -1988
rect 13026 -2090 13060 -2056
rect 13026 -2158 13060 -2124
rect 13026 -2226 13060 -2192
rect 13026 -2294 13060 -2260
rect 13026 -2362 13060 -2328
rect 13026 -2430 13060 -2396
rect 13026 -2498 13060 -2464
rect 13026 -2566 13060 -2532
rect 13026 -2634 13060 -2600
rect 13026 -2702 13060 -2668
rect 13026 -2770 13060 -2736
rect 13026 -2838 13060 -2804
rect 13026 -2906 13060 -2872
rect 13430 -2022 13464 -1988
rect 13430 -2090 13464 -2056
rect 13430 -2158 13464 -2124
rect 13430 -2226 13464 -2192
rect 13430 -2294 13464 -2260
rect 13430 -2362 13464 -2328
rect 13430 -2430 13464 -2396
rect 13430 -2498 13464 -2464
rect 13430 -2566 13464 -2532
rect 13430 -2634 13464 -2600
rect 13430 -2702 13464 -2668
rect 13430 -2770 13464 -2736
rect 13430 -2838 13464 -2804
rect 13430 -2906 13464 -2872
<< poly >>
rect 11380 -3414 11410 -3348
rect 11716 -3414 11746 -3348
rect 12052 -3414 12082 -3348
rect 12388 -3414 12418 -3348
rect 12724 -3414 12754 -3348
rect 13060 -3414 13090 -3348
<< locali >>
rect 11006 -1972 11040 -1956
rect 11006 -2964 11040 -2948
rect 11410 -1972 11444 -1956
rect 11410 -2964 11444 -2948
rect 11814 -1972 11848 -1956
rect 11814 -2964 11848 -2948
rect 12218 -1972 12252 -1956
rect 12218 -2964 12252 -2948
rect 12622 -1972 12656 -1956
rect 12622 -2964 12656 -2948
rect 13026 -1972 13060 -1956
rect 13026 -2964 13060 -2948
rect 13430 -1972 13464 -1956
rect 13430 -2964 13464 -2948
rect 11380 -3398 11410 -3364
rect 11716 -3398 11746 -3364
rect 12052 -3398 12082 -3364
rect 12388 -3398 12418 -3364
rect 12724 -3398 12754 -3364
rect 13060 -3398 13090 -3364
rect 11210 -3490 11244 -3432
rect 11210 -3558 11244 -3524
rect 11210 -3626 11244 -3592
rect 11210 -3694 11244 -3660
rect 11210 -3736 11244 -3728
rect 11210 -4440 11244 -4424
rect 11546 -3464 11580 -3432
rect 11546 -3532 11580 -3498
rect 11546 -3600 11580 -3566
rect 11546 -3668 11580 -3634
rect 11546 -3736 11580 -3702
rect 11546 -4440 11580 -4424
rect 11882 -3464 11916 -3432
rect 11882 -3532 11916 -3498
rect 11882 -3600 11916 -3566
rect 11882 -3668 11916 -3634
rect 11882 -3736 11916 -3702
rect 11882 -4440 11916 -4424
rect 12218 -3464 12252 -3432
rect 12218 -3532 12252 -3498
rect 12218 -3600 12252 -3566
rect 12218 -3668 12252 -3634
rect 12218 -3736 12252 -3702
rect 12218 -4440 12252 -4424
rect 12554 -3464 12588 -3432
rect 12554 -3532 12588 -3498
rect 12554 -3600 12588 -3566
rect 12554 -3668 12588 -3634
rect 12554 -3736 12588 -3702
rect 12554 -4440 12588 -4424
rect 12890 -3464 12924 -3432
rect 12890 -3532 12924 -3498
rect 12890 -3600 12924 -3566
rect 12890 -3668 12924 -3634
rect 12890 -3736 12924 -3702
rect 12890 -4440 12924 -4424
rect 13226 -3464 13260 -3432
rect 13226 -3532 13260 -3498
rect 13226 -3600 13260 -3566
rect 13226 -3668 13260 -3634
rect 13226 -3736 13260 -3702
rect 13226 -4440 13260 -4424
<< viali >>
rect 11006 -2014 11040 -1972
rect 11006 -2048 11040 -2014
rect 11006 -2082 11040 -2048
rect 11006 -2116 11040 -2082
rect 11006 -2150 11040 -2116
rect 11006 -2184 11040 -2150
rect 11006 -2218 11040 -2184
rect 11006 -2252 11040 -2218
rect 11006 -2286 11040 -2252
rect 11006 -2320 11040 -2286
rect 11006 -2354 11040 -2320
rect 11006 -2388 11040 -2354
rect 11006 -2422 11040 -2388
rect 11006 -2456 11040 -2422
rect 11006 -2490 11040 -2456
rect 11006 -2524 11040 -2490
rect 11006 -2558 11040 -2524
rect 11006 -2592 11040 -2558
rect 11006 -2626 11040 -2592
rect 11006 -2660 11040 -2626
rect 11006 -2694 11040 -2660
rect 11006 -2728 11040 -2694
rect 11006 -2762 11040 -2728
rect 11006 -2796 11040 -2762
rect 11006 -2830 11040 -2796
rect 11006 -2864 11040 -2830
rect 11006 -2898 11040 -2864
rect 11006 -2932 11040 -2898
rect 11006 -2948 11040 -2932
rect 11410 -1988 11444 -1972
rect 11410 -2022 11444 -1988
rect 11410 -2056 11444 -2022
rect 11410 -2090 11444 -2056
rect 11410 -2124 11444 -2090
rect 11410 -2158 11444 -2124
rect 11410 -2192 11444 -2158
rect 11410 -2226 11444 -2192
rect 11410 -2260 11444 -2226
rect 11410 -2294 11444 -2260
rect 11410 -2328 11444 -2294
rect 11410 -2362 11444 -2328
rect 11410 -2396 11444 -2362
rect 11410 -2430 11444 -2396
rect 11410 -2464 11444 -2430
rect 11410 -2498 11444 -2464
rect 11410 -2532 11444 -2498
rect 11410 -2566 11444 -2532
rect 11410 -2600 11444 -2566
rect 11410 -2634 11444 -2600
rect 11410 -2668 11444 -2634
rect 11410 -2702 11444 -2668
rect 11410 -2736 11444 -2702
rect 11410 -2770 11444 -2736
rect 11410 -2804 11444 -2770
rect 11410 -2838 11444 -2804
rect 11410 -2872 11444 -2838
rect 11410 -2906 11444 -2872
rect 11410 -2948 11444 -2906
rect 11814 -1988 11848 -1972
rect 11814 -2022 11848 -1988
rect 11814 -2056 11848 -2022
rect 11814 -2090 11848 -2056
rect 11814 -2124 11848 -2090
rect 11814 -2158 11848 -2124
rect 11814 -2192 11848 -2158
rect 11814 -2226 11848 -2192
rect 11814 -2260 11848 -2226
rect 11814 -2294 11848 -2260
rect 11814 -2328 11848 -2294
rect 11814 -2362 11848 -2328
rect 11814 -2396 11848 -2362
rect 11814 -2430 11848 -2396
rect 11814 -2464 11848 -2430
rect 11814 -2498 11848 -2464
rect 11814 -2532 11848 -2498
rect 11814 -2566 11848 -2532
rect 11814 -2600 11848 -2566
rect 11814 -2634 11848 -2600
rect 11814 -2668 11848 -2634
rect 11814 -2702 11848 -2668
rect 11814 -2736 11848 -2702
rect 11814 -2770 11848 -2736
rect 11814 -2804 11848 -2770
rect 11814 -2838 11848 -2804
rect 11814 -2872 11848 -2838
rect 11814 -2906 11848 -2872
rect 11814 -2948 11848 -2906
rect 12218 -1988 12252 -1972
rect 12218 -2022 12252 -1988
rect 12218 -2056 12252 -2022
rect 12218 -2090 12252 -2056
rect 12218 -2124 12252 -2090
rect 12218 -2158 12252 -2124
rect 12218 -2192 12252 -2158
rect 12218 -2226 12252 -2192
rect 12218 -2260 12252 -2226
rect 12218 -2294 12252 -2260
rect 12218 -2328 12252 -2294
rect 12218 -2362 12252 -2328
rect 12218 -2396 12252 -2362
rect 12218 -2430 12252 -2396
rect 12218 -2464 12252 -2430
rect 12218 -2498 12252 -2464
rect 12218 -2532 12252 -2498
rect 12218 -2566 12252 -2532
rect 12218 -2600 12252 -2566
rect 12218 -2634 12252 -2600
rect 12218 -2668 12252 -2634
rect 12218 -2702 12252 -2668
rect 12218 -2736 12252 -2702
rect 12218 -2770 12252 -2736
rect 12218 -2804 12252 -2770
rect 12218 -2838 12252 -2804
rect 12218 -2872 12252 -2838
rect 12218 -2906 12252 -2872
rect 12218 -2948 12252 -2906
rect 12622 -1988 12656 -1972
rect 12622 -2022 12656 -1988
rect 12622 -2056 12656 -2022
rect 12622 -2090 12656 -2056
rect 12622 -2124 12656 -2090
rect 12622 -2158 12656 -2124
rect 12622 -2192 12656 -2158
rect 12622 -2226 12656 -2192
rect 12622 -2260 12656 -2226
rect 12622 -2294 12656 -2260
rect 12622 -2328 12656 -2294
rect 12622 -2362 12656 -2328
rect 12622 -2396 12656 -2362
rect 12622 -2430 12656 -2396
rect 12622 -2464 12656 -2430
rect 12622 -2498 12656 -2464
rect 12622 -2532 12656 -2498
rect 12622 -2566 12656 -2532
rect 12622 -2600 12656 -2566
rect 12622 -2634 12656 -2600
rect 12622 -2668 12656 -2634
rect 12622 -2702 12656 -2668
rect 12622 -2736 12656 -2702
rect 12622 -2770 12656 -2736
rect 12622 -2804 12656 -2770
rect 12622 -2838 12656 -2804
rect 12622 -2872 12656 -2838
rect 12622 -2906 12656 -2872
rect 12622 -2948 12656 -2906
rect 13026 -1988 13060 -1972
rect 13026 -2022 13060 -1988
rect 13026 -2056 13060 -2022
rect 13026 -2090 13060 -2056
rect 13026 -2124 13060 -2090
rect 13026 -2158 13060 -2124
rect 13026 -2192 13060 -2158
rect 13026 -2226 13060 -2192
rect 13026 -2260 13060 -2226
rect 13026 -2294 13060 -2260
rect 13026 -2328 13060 -2294
rect 13026 -2362 13060 -2328
rect 13026 -2396 13060 -2362
rect 13026 -2430 13060 -2396
rect 13026 -2464 13060 -2430
rect 13026 -2498 13060 -2464
rect 13026 -2532 13060 -2498
rect 13026 -2566 13060 -2532
rect 13026 -2600 13060 -2566
rect 13026 -2634 13060 -2600
rect 13026 -2668 13060 -2634
rect 13026 -2702 13060 -2668
rect 13026 -2736 13060 -2702
rect 13026 -2770 13060 -2736
rect 13026 -2804 13060 -2770
rect 13026 -2838 13060 -2804
rect 13026 -2872 13060 -2838
rect 13026 -2906 13060 -2872
rect 13026 -2948 13060 -2906
rect 13430 -1988 13464 -1972
rect 13430 -2022 13464 -1988
rect 13430 -2056 13464 -2022
rect 13430 -2090 13464 -2056
rect 13430 -2124 13464 -2090
rect 13430 -2158 13464 -2124
rect 13430 -2192 13464 -2158
rect 13430 -2226 13464 -2192
rect 13430 -2260 13464 -2226
rect 13430 -2294 13464 -2260
rect 13430 -2328 13464 -2294
rect 13430 -2362 13464 -2328
rect 13430 -2396 13464 -2362
rect 13430 -2430 13464 -2396
rect 13430 -2464 13464 -2430
rect 13430 -2498 13464 -2464
rect 13430 -2532 13464 -2498
rect 13430 -2566 13464 -2532
rect 13430 -2600 13464 -2566
rect 13430 -2634 13464 -2600
rect 13430 -2668 13464 -2634
rect 13430 -2702 13464 -2668
rect 13430 -2736 13464 -2702
rect 13430 -2770 13464 -2736
rect 13430 -2804 13464 -2770
rect 13430 -2838 13464 -2804
rect 13430 -2872 13464 -2838
rect 13430 -2906 13464 -2872
rect 13430 -2948 13464 -2906
rect 11210 -3762 11244 -3736
rect 11210 -3796 11244 -3762
rect 11210 -3830 11244 -3796
rect 11210 -3864 11244 -3830
rect 11210 -3898 11244 -3864
rect 11210 -3932 11244 -3898
rect 11210 -3966 11244 -3932
rect 11210 -4000 11244 -3966
rect 11210 -4034 11244 -4000
rect 11210 -4068 11244 -4034
rect 11210 -4102 11244 -4068
rect 11210 -4136 11244 -4102
rect 11210 -4170 11244 -4136
rect 11210 -4204 11244 -4170
rect 11210 -4238 11244 -4204
rect 11210 -4272 11244 -4238
rect 11210 -4306 11244 -4272
rect 11210 -4340 11244 -4306
rect 11210 -4374 11244 -4340
rect 11210 -4408 11244 -4374
rect 11210 -4424 11244 -4408
rect 11546 -3770 11580 -3736
rect 11546 -3804 11580 -3770
rect 11546 -3838 11580 -3804
rect 11546 -3872 11580 -3838
rect 11546 -3906 11580 -3872
rect 11546 -3940 11580 -3906
rect 11546 -3974 11580 -3940
rect 11546 -4008 11580 -3974
rect 11546 -4042 11580 -4008
rect 11546 -4076 11580 -4042
rect 11546 -4110 11580 -4076
rect 11546 -4144 11580 -4110
rect 11546 -4178 11580 -4144
rect 11546 -4212 11580 -4178
rect 11546 -4246 11580 -4212
rect 11546 -4280 11580 -4246
rect 11546 -4314 11580 -4280
rect 11546 -4348 11580 -4314
rect 11546 -4382 11580 -4348
rect 11546 -4424 11580 -4382
rect 11882 -3770 11916 -3736
rect 11882 -3804 11916 -3770
rect 11882 -3838 11916 -3804
rect 11882 -3872 11916 -3838
rect 11882 -3906 11916 -3872
rect 11882 -3940 11916 -3906
rect 11882 -3974 11916 -3940
rect 11882 -4008 11916 -3974
rect 11882 -4042 11916 -4008
rect 11882 -4076 11916 -4042
rect 11882 -4110 11916 -4076
rect 11882 -4144 11916 -4110
rect 11882 -4178 11916 -4144
rect 11882 -4212 11916 -4178
rect 11882 -4246 11916 -4212
rect 11882 -4280 11916 -4246
rect 11882 -4314 11916 -4280
rect 11882 -4348 11916 -4314
rect 11882 -4382 11916 -4348
rect 11882 -4424 11916 -4382
rect 12218 -3770 12252 -3736
rect 12218 -3804 12252 -3770
rect 12218 -3838 12252 -3804
rect 12218 -3872 12252 -3838
rect 12218 -3906 12252 -3872
rect 12218 -3940 12252 -3906
rect 12218 -3974 12252 -3940
rect 12218 -4008 12252 -3974
rect 12218 -4042 12252 -4008
rect 12218 -4076 12252 -4042
rect 12218 -4110 12252 -4076
rect 12218 -4144 12252 -4110
rect 12218 -4178 12252 -4144
rect 12218 -4212 12252 -4178
rect 12218 -4246 12252 -4212
rect 12218 -4280 12252 -4246
rect 12218 -4314 12252 -4280
rect 12218 -4348 12252 -4314
rect 12218 -4382 12252 -4348
rect 12218 -4424 12252 -4382
rect 12554 -3770 12588 -3736
rect 12554 -3804 12588 -3770
rect 12554 -3838 12588 -3804
rect 12554 -3872 12588 -3838
rect 12554 -3906 12588 -3872
rect 12554 -3940 12588 -3906
rect 12554 -3974 12588 -3940
rect 12554 -4008 12588 -3974
rect 12554 -4042 12588 -4008
rect 12554 -4076 12588 -4042
rect 12554 -4110 12588 -4076
rect 12554 -4144 12588 -4110
rect 12554 -4178 12588 -4144
rect 12554 -4212 12588 -4178
rect 12554 -4246 12588 -4212
rect 12554 -4280 12588 -4246
rect 12554 -4314 12588 -4280
rect 12554 -4348 12588 -4314
rect 12554 -4382 12588 -4348
rect 12554 -4424 12588 -4382
rect 12890 -3770 12924 -3736
rect 12890 -3804 12924 -3770
rect 12890 -3838 12924 -3804
rect 12890 -3872 12924 -3838
rect 12890 -3906 12924 -3872
rect 12890 -3940 12924 -3906
rect 12890 -3974 12924 -3940
rect 12890 -4008 12924 -3974
rect 12890 -4042 12924 -4008
rect 12890 -4076 12924 -4042
rect 12890 -4110 12924 -4076
rect 12890 -4144 12924 -4110
rect 12890 -4178 12924 -4144
rect 12890 -4212 12924 -4178
rect 12890 -4246 12924 -4212
rect 12890 -4280 12924 -4246
rect 12890 -4314 12924 -4280
rect 12890 -4348 12924 -4314
rect 12890 -4382 12924 -4348
rect 12890 -4424 12924 -4382
rect 13226 -3770 13260 -3736
rect 13226 -3804 13260 -3770
rect 13226 -3838 13260 -3804
rect 13226 -3872 13260 -3838
rect 13226 -3906 13260 -3872
rect 13226 -3940 13260 -3906
rect 13226 -3974 13260 -3940
rect 13226 -4008 13260 -3974
rect 13226 -4042 13260 -4008
rect 13226 -4076 13260 -4042
rect 13226 -4110 13260 -4076
rect 13226 -4144 13260 -4110
rect 13226 -4178 13260 -4144
rect 13226 -4212 13260 -4178
rect 13226 -4246 13260 -4212
rect 13226 -4280 13260 -4246
rect 13226 -4314 13260 -4280
rect 13226 -4348 13260 -4314
rect 13226 -4382 13260 -4348
rect 13226 -4424 13260 -4382
<< metal1 >>
rect 10846 -1498 10958 -1488
rect 10846 -1666 10876 -1498
rect 10932 -1666 10958 -1498
rect 10846 -3248 10958 -1666
rect 10986 -1768 13482 -1762
rect 10986 -1820 11006 -1768
rect 13462 -1820 13482 -1768
rect 10986 -1826 13482 -1820
rect 10986 -1972 11098 -1826
rect 10986 -2948 11006 -1972
rect 11040 -2948 11098 -1972
rect 10986 -2960 11098 -2948
rect 11196 -1972 11254 -1962
rect 11196 -2954 11254 -2948
rect 11370 -1972 11482 -1826
rect 11370 -2948 11410 -1972
rect 11444 -2948 11482 -1972
rect 11370 -2960 11482 -2948
rect 11600 -1972 11658 -1962
rect 11600 -2954 11658 -2948
rect 11774 -1972 11886 -1826
rect 11774 -2948 11814 -1972
rect 11848 -2948 11886 -1972
rect 11774 -2960 11886 -2948
rect 12004 -1972 12062 -1962
rect 12004 -2954 12062 -2948
rect 12178 -1972 12290 -1826
rect 12178 -2948 12218 -1972
rect 12252 -2948 12290 -1972
rect 12178 -2960 12290 -2948
rect 12408 -1972 12466 -1962
rect 12408 -2954 12466 -2948
rect 12582 -1972 12694 -1826
rect 12582 -2948 12622 -1972
rect 12656 -2948 12694 -1972
rect 12582 -2960 12694 -2948
rect 12812 -1972 12870 -1962
rect 12812 -2954 12870 -2948
rect 12986 -1972 13098 -1826
rect 12986 -2948 13026 -1972
rect 13060 -2948 13098 -1972
rect 12986 -2960 13098 -2948
rect 13216 -1972 13274 -1962
rect 13216 -2954 13274 -2948
rect 13370 -1972 13482 -1826
rect 13370 -2948 13430 -1972
rect 13464 -2948 13482 -1972
rect 13370 -2960 13482 -2948
rect 11128 -3060 11322 -3000
rect 11532 -3060 11726 -3000
rect 11200 -3102 11322 -3060
rect 11200 -3108 11450 -3102
rect 11424 -3160 11450 -3108
rect 11200 -3166 11450 -3160
rect 10846 -3306 10958 -3300
rect 11316 -3348 11450 -3166
rect 11562 -3242 11696 -3060
rect 11936 -3102 12130 -3000
rect 11936 -3108 12160 -3102
rect 11936 -3166 12160 -3160
rect 11562 -3248 11810 -3242
rect 11786 -3300 11810 -3248
rect 11562 -3306 11810 -3300
rect 11316 -3404 11474 -3348
rect 11652 -3404 11810 -3306
rect 11988 -3404 12146 -3166
rect 12340 -3242 12534 -3000
rect 12744 -3102 12938 -3000
rect 12690 -3108 12938 -3102
rect 12914 -3160 12938 -3108
rect 12690 -3166 12938 -3160
rect 13148 -3078 13342 -3000
rect 12316 -3248 12540 -3242
rect 12316 -3306 12540 -3300
rect 12324 -3404 12482 -3306
rect 12690 -3348 12802 -3166
rect 13148 -3242 13268 -3078
rect 13036 -3248 13268 -3242
rect 13260 -3300 13268 -3248
rect 13036 -3306 13268 -3300
rect 13376 -3108 13488 -3102
rect 13036 -3348 13154 -3306
rect 12660 -3404 12818 -3348
rect 12996 -3404 13154 -3348
rect 8712 -4564 9216 -3706
rect 11188 -3728 11244 -3436
rect 11272 -3442 11330 -3436
rect 11272 -3706 11330 -3700
rect 11460 -3442 11518 -3436
rect 11460 -3706 11518 -3700
rect 11188 -3736 11250 -3728
rect 11546 -3730 11580 -3436
rect 11608 -3442 11666 -3436
rect 11608 -3706 11666 -3700
rect 11796 -3442 11854 -3436
rect 11796 -3706 11854 -3700
rect 11882 -3730 11916 -3436
rect 11944 -3442 12002 -3436
rect 11944 -3706 12002 -3700
rect 12132 -3442 12190 -3436
rect 12132 -3706 12190 -3700
rect 12218 -3730 12252 -3436
rect 12280 -3442 12338 -3436
rect 12280 -3706 12338 -3700
rect 12468 -3442 12526 -3436
rect 12468 -3706 12526 -3700
rect 12554 -3730 12588 -3436
rect 12616 -3442 12674 -3436
rect 12616 -3706 12674 -3700
rect 12804 -3442 12862 -3436
rect 12804 -3706 12862 -3700
rect 12890 -3730 12924 -3436
rect 12952 -3442 13010 -3436
rect 12952 -3706 13010 -3700
rect 13140 -3442 13198 -3436
rect 13140 -3706 13198 -3700
rect 13226 -3730 13282 -3436
rect 11188 -4424 11210 -3736
rect 11244 -4424 11250 -3736
rect 11540 -3736 11586 -3730
rect 11188 -4558 11250 -4424
rect 11366 -4050 11424 -4040
rect 11366 -4436 11424 -4422
rect 11540 -4424 11546 -3736
rect 11580 -4424 11586 -3736
rect 11876 -3736 11922 -3730
rect 11540 -4558 11586 -4424
rect 11702 -4050 11760 -4040
rect 11702 -4436 11760 -4422
rect 11876 -4424 11882 -3736
rect 11916 -4424 11922 -3736
rect 12212 -3736 12258 -3730
rect 11876 -4558 11922 -4424
rect 12038 -4050 12096 -4040
rect 12038 -4436 12096 -4422
rect 12212 -4424 12218 -3736
rect 12252 -4424 12258 -3736
rect 12548 -3736 12594 -3730
rect 12212 -4558 12258 -4424
rect 12374 -4050 12432 -4040
rect 12374 -4436 12432 -4422
rect 12548 -4424 12554 -3736
rect 12588 -4424 12594 -3736
rect 12884 -3736 12930 -3730
rect 12548 -4558 12594 -4424
rect 12710 -4050 12768 -4040
rect 12710 -4436 12768 -4422
rect 12884 -4424 12890 -3736
rect 12924 -4424 12930 -3736
rect 13220 -3736 13282 -3730
rect 12884 -4558 12930 -4424
rect 13046 -4050 13104 -4040
rect 13046 -4436 13104 -4422
rect 13220 -4424 13226 -3736
rect 13260 -4424 13282 -3736
rect 13220 -4558 13282 -4424
rect 8712 -4616 8740 -4564
rect 9188 -4616 9216 -4564
rect 8712 -4646 9216 -4616
rect 11172 -4564 13296 -4558
rect 11172 -4616 11192 -4564
rect 13276 -4616 13296 -4564
rect 11172 -4622 13296 -4616
rect 13376 -4708 13488 -3160
rect 13376 -4876 13404 -4708
rect 13460 -4876 13488 -4708
rect 13376 -4886 13488 -4876
<< via1 >>
rect 10876 -1666 10932 -1498
rect 11006 -1820 13462 -1768
rect 11196 -2948 11254 -1972
rect 11600 -2948 11658 -1972
rect 12004 -2948 12062 -1972
rect 12408 -2948 12466 -1972
rect 12812 -2948 12870 -1972
rect 13216 -2948 13274 -1972
rect 11200 -3160 11424 -3108
rect 10846 -3300 10958 -3248
rect 11936 -3160 12160 -3108
rect 11562 -3300 11786 -3248
rect 12690 -3160 12914 -3108
rect 12316 -3300 12540 -3248
rect 13036 -3300 13260 -3248
rect 13376 -3160 13488 -3108
rect 11272 -3700 11330 -3442
rect 11460 -3700 11518 -3442
rect 11608 -3700 11666 -3442
rect 11796 -3700 11854 -3442
rect 11944 -3700 12002 -3442
rect 12132 -3700 12190 -3442
rect 12280 -3700 12338 -3442
rect 12468 -3700 12526 -3442
rect 12616 -3700 12674 -3442
rect 12804 -3700 12862 -3442
rect 12952 -3700 13010 -3442
rect 13140 -3700 13198 -3442
rect 11366 -4422 11424 -4050
rect 11702 -4422 11760 -4050
rect 12038 -4422 12096 -4050
rect 12374 -4422 12432 -4050
rect 12710 -4422 12768 -4050
rect 13046 -4422 13104 -4050
rect 8740 -4616 9188 -4564
rect 11192 -4616 13276 -4564
rect 13404 -4876 13460 -4708
<< metal2 >>
rect 10846 -1498 10958 -1488
rect 10846 -1666 10876 -1498
rect 10932 -1666 10958 -1498
rect 10846 -1676 10958 -1666
rect 10986 -1768 14160 -1710
rect 10986 -1820 11006 -1768
rect 13462 -1774 14160 -1768
rect 13462 -1790 14136 -1774
rect 13462 -1820 13968 -1790
rect 10986 -1878 13968 -1820
rect 11196 -1972 11254 -1962
rect 11196 -2960 11254 -2948
rect 11600 -1972 11658 -1962
rect 11600 -2960 11658 -2948
rect 12004 -1972 12062 -1962
rect 12004 -2960 12062 -2948
rect 12408 -1972 12466 -1962
rect 12408 -2960 12466 -2948
rect 12812 -1972 12870 -1962
rect 12812 -2960 12870 -2948
rect 13216 -1972 13274 -1962
rect 13216 -2960 13274 -2948
rect 11200 -3078 11322 -3050
rect 11122 -3108 13488 -3078
rect 11122 -3160 11200 -3108
rect 11424 -3160 11936 -3108
rect 12160 -3160 12690 -3108
rect 12914 -3160 13376 -3108
rect 11122 -3190 13488 -3160
rect 10846 -3248 13348 -3218
rect 10958 -3300 11562 -3248
rect 11786 -3300 12316 -3248
rect 12540 -3300 13036 -3248
rect 13260 -3300 13348 -3248
rect 10846 -3330 13348 -3300
rect 8712 -3442 13198 -3436
rect 8712 -3486 11272 -3442
rect 8712 -3598 8756 -3486
rect 9750 -3598 11272 -3486
rect 8712 -3660 11272 -3598
rect 11330 -3660 11460 -3442
rect 11272 -3706 11330 -3700
rect 11518 -3660 11608 -3442
rect 11460 -3706 11518 -3700
rect 11666 -3660 11796 -3442
rect 11608 -3706 11666 -3700
rect 11854 -3660 11944 -3442
rect 11796 -3706 11854 -3700
rect 12002 -3660 12132 -3442
rect 11944 -3706 12002 -3700
rect 12190 -3660 12280 -3442
rect 12132 -3706 12190 -3700
rect 12338 -3660 12468 -3442
rect 12280 -3706 12338 -3700
rect 12526 -3660 12616 -3442
rect 12468 -3706 12526 -3700
rect 12674 -3660 12804 -3442
rect 12616 -3706 12674 -3700
rect 12862 -3660 12952 -3442
rect 12804 -3706 12862 -3700
rect 13010 -3660 13140 -3442
rect 12952 -3706 13010 -3700
rect 13140 -3706 13198 -3700
rect 13912 -3758 13968 -1878
rect 14080 -3758 14136 -1790
rect 13912 -3774 14136 -3758
rect 11366 -4050 11424 -4040
rect 11366 -4436 11424 -4422
rect 11702 -4050 11760 -4040
rect 11702 -4436 11760 -4422
rect 12038 -4050 12096 -4040
rect 12038 -4436 12096 -4422
rect 12374 -4050 12432 -4040
rect 12374 -4436 12432 -4422
rect 12710 -4050 12768 -4040
rect 12710 -4436 12768 -4422
rect 13046 -4050 13104 -4040
rect 13046 -4436 13104 -4422
rect 8712 -4564 13296 -4534
rect 8712 -4616 8740 -4564
rect 9188 -4616 11192 -4564
rect 13276 -4616 13296 -4564
rect 8712 -4646 13296 -4616
rect 13376 -4708 13488 -4698
rect 13376 -4876 13404 -4708
rect 13460 -4876 13488 -4708
rect 13376 -4886 13488 -4876
<< via2 >>
rect 10876 -1666 10932 -1498
rect 11196 -2948 11254 -1972
rect 11600 -2948 11658 -1972
rect 12004 -2948 12062 -1972
rect 12408 -2948 12466 -1972
rect 12812 -2948 12870 -1972
rect 13216 -2948 13274 -1972
rect 8756 -3598 9750 -3486
rect 13968 -3758 14080 -1790
rect 11366 -4422 11424 -4050
rect 11702 -4422 11760 -4050
rect 12038 -4422 12096 -4050
rect 12374 -4422 12432 -4050
rect 12710 -4422 12768 -4050
rect 13046 -4422 13104 -4050
rect 13404 -4876 13460 -4708
<< metal3 >>
rect 8812 -1498 14892 -1454
rect 8812 -1666 10876 -1498
rect 10932 -1666 14892 -1498
rect 8812 -1694 14892 -1666
rect 8712 -3486 9792 -1774
rect 8712 -3598 8756 -3486
rect 9750 -3598 9792 -3486
rect 8712 -3660 9792 -3598
rect 11190 -1972 11370 -1694
rect 11190 -2948 11196 -1972
rect 11254 -2948 11370 -1972
rect 11190 -3440 11370 -2948
rect 11594 -1972 11774 -1960
rect 11594 -2948 11600 -1972
rect 11658 -2948 11774 -1972
rect 11190 -4050 11430 -3440
rect 11190 -4422 11366 -4050
rect 11424 -4422 11430 -4050
rect 11190 -4428 11430 -4422
rect 11594 -4050 11774 -2948
rect 11594 -4422 11702 -4050
rect 11760 -4422 11774 -4050
rect 11594 -4682 11774 -4422
rect 11998 -1972 12178 -1694
rect 11998 -2948 12004 -1972
rect 12062 -2948 12178 -1972
rect 11998 -4050 12178 -2948
rect 11998 -4422 12038 -4050
rect 12096 -4422 12178 -4050
rect 11998 -4428 12178 -4422
rect 12352 -1972 12532 -1960
rect 12352 -2948 12408 -1972
rect 12466 -2948 12532 -1972
rect 12352 -4050 12532 -2948
rect 12352 -4422 12374 -4050
rect 12432 -4422 12532 -4050
rect 12352 -4682 12532 -4422
rect 12696 -1972 12876 -1694
rect 13912 -1790 14992 -1774
rect 12696 -2948 12812 -1972
rect 12870 -2948 12876 -1972
rect 12696 -4050 12876 -2948
rect 12696 -4422 12710 -4050
rect 12768 -4422 12876 -4050
rect 12696 -4428 12876 -4422
rect 13040 -1972 13280 -1960
rect 13040 -2948 13216 -1972
rect 13274 -2948 13280 -1972
rect 13040 -2960 13280 -2948
rect 13040 -4050 13226 -2960
rect 13912 -3758 13968 -1790
rect 14080 -3758 14992 -1790
rect 13912 -3774 14992 -3758
rect 13040 -4422 13046 -4050
rect 13104 -4422 13226 -4050
rect 13040 -4682 13226 -4422
rect 8812 -4708 14892 -4682
rect 8812 -4766 13404 -4708
rect 13460 -4766 14892 -4708
rect 8812 -4836 8818 -4766
rect 14882 -4836 14892 -4766
rect 8812 -4876 13404 -4836
rect 13460 -4876 14892 -4836
rect 8812 -4922 14892 -4876
<< via3 >>
rect 8818 -4836 13404 -4766
rect 13404 -4836 13460 -4766
rect 13460 -4836 14882 -4766
<< metal4 >>
rect 8712 4928 14992 6008
rect 8892 4816 14812 4928
rect 8812 -4766 14892 -4760
rect 8812 -4836 8818 -4766
rect 14882 -4836 14892 -4766
rect 8812 -5086 14892 -4836
rect 8712 -11394 14994 -11280
rect 8712 -12474 14992 -11394
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M11
timestamp 1681062556
transform 1 0 11348 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M12
timestamp 1681062556
transform 1 0 11442 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M13
timestamp 1681062556
transform 1 0 12020 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M14
timestamp 1681062556
transform 1 0 12114 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M15
timestamp 1681062556
transform 1 0 12692 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M16
timestamp 1681062556
transform 1 0 12786 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M21
timestamp 1681062556
transform 1 0 11684 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M22
timestamp 1681062556
transform 1 0 11778 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M23
timestamp 1681062556
transform 1 0 12356 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M24
timestamp 1681062556
transform 1 0 12450 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M25
timestamp 1681062556
transform 1 0 13028 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__nfet_01v8_lvt_R7ME6Q  M26
timestamp 1681062556
transform 1 0 13122 0 1 -3905
box -76 -557 76 557
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M31
timestamp 1681050310
transform 1 0 11161 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M32
timestamp 1681050310
transform 1 0 11289 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M33
timestamp 1681050310
transform 1 0 11969 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M34
timestamp 1681050310
transform 1 0 12097 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M35
timestamp 1681050310
transform 1 0 12777 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M36
timestamp 1681050310
transform 1 0 12905 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M41
timestamp 1681050310
transform 1 0 11565 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M42
timestamp 1681050310
transform 1 0 11693 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M43
timestamp 1681050310
transform 1 0 12373 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M44
timestamp 1681050310
transform 1 0 12501 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M45
timestamp 1681050310
transform 1 0 13181 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__pfet_01v8_lvt_73FV24  M46
timestamp 1681050310
transform 1 0 13309 0 1 -2496
box -129 -564 129 598
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1680390383
transform 0 1 11852 -1 0 1722
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 1680390383
transform 0 1 11852 -1 0 -8188
box -3186 -3040 3186 3040
<< labels >>
flabel metal1 8712 -4646 9216 -3706 0 FreeMono 1280 0 0 0 vss
port 4 nsew
flabel metal3 8712 -3660 9792 -1774 0 FreeMono 1920 0 0 0 out1
port 2 nsew
flabel metal3 13912 -3774 14992 -1774 0 FreeMono 1920 0 0 0 out2
port 3 nsew
flabel metal4 8712 4928 14992 6008 0 FreeMono 3200 0 0 0 vinp
port 0 nsew
flabel metal4 8712 -12474 14992 -11394 0 FreeMono 3200 0 0 0 vinn
port 1 nsew
<< end >>
