magic
tech sky130A
magscale 1 2
timestamp 1681766136
<< nwell >>
rect 3918 -576 3984 586
rect 4982 -576 5096 586
rect 5634 -576 5700 586
rect 6698 -576 6812 586
rect 7810 -576 7876 586
rect 3918 -2446 3984 -1284
rect 4982 -2446 5096 -1284
rect 5636 -2446 5702 -1284
rect 6700 -2446 6814 -1284
rect 7812 -2446 7878 -1284
<< ndiff >>
rect 3608 -3426 3610 -3026
rect 4584 -3426 4586 -3026
rect 4672 -3426 4674 -3026
rect 5648 -3426 5650 -3026
rect 5736 -3426 5738 -3026
rect 6712 -3426 6714 -3026
rect 6800 -3426 6802 -3026
rect 7776 -3426 7778 -3026
rect 7864 -3426 7866 -3026
<< pdiff >>
rect 4018 -476 4020 524
rect 4994 -476 4996 524
rect 5082 -476 5084 524
rect 5734 -476 5736 524
rect 6710 -476 6712 524
rect 6798 -476 6800 524
rect 7774 -476 7776 524
rect 4018 -2384 4020 -1384
rect 4994 -2384 4996 -1384
rect 5082 -2384 5084 -1384
rect 5736 -2384 5738 -1384
rect 6712 -2384 6714 -1384
rect 6800 -2384 6802 -1384
rect 7776 -2384 7778 -1384
<< psubdiff >>
rect 3544 -3092 3608 -3026
rect 3544 -3126 3548 -3092
rect 3582 -3126 3608 -3092
rect 3544 -3160 3608 -3126
rect 3544 -3194 3548 -3160
rect 3582 -3194 3608 -3160
rect 3544 -3228 3608 -3194
rect 3544 -3262 3548 -3228
rect 3582 -3262 3608 -3228
rect 3544 -3296 3608 -3262
rect 3544 -3330 3548 -3296
rect 3582 -3330 3608 -3296
rect 3544 -3364 3608 -3330
rect 3544 -3398 3548 -3364
rect 3582 -3398 3608 -3364
rect 3544 -3426 3608 -3398
rect 4586 -3092 4672 -3026
rect 4586 -3126 4612 -3092
rect 4646 -3126 4672 -3092
rect 4586 -3160 4672 -3126
rect 4586 -3194 4612 -3160
rect 4646 -3194 4672 -3160
rect 4586 -3228 4672 -3194
rect 4586 -3262 4612 -3228
rect 4646 -3262 4672 -3228
rect 4586 -3296 4672 -3262
rect 4586 -3330 4612 -3296
rect 4646 -3330 4672 -3296
rect 4586 -3364 4672 -3330
rect 4586 -3398 4612 -3364
rect 4646 -3398 4672 -3364
rect 4586 -3426 4672 -3398
rect 5650 -3092 5736 -3026
rect 5650 -3126 5676 -3092
rect 5710 -3126 5736 -3092
rect 5650 -3160 5736 -3126
rect 5650 -3194 5676 -3160
rect 5710 -3194 5736 -3160
rect 5650 -3228 5736 -3194
rect 5650 -3262 5676 -3228
rect 5710 -3262 5736 -3228
rect 5650 -3296 5736 -3262
rect 5650 -3330 5676 -3296
rect 5710 -3330 5736 -3296
rect 5650 -3364 5736 -3330
rect 5650 -3398 5676 -3364
rect 5710 -3398 5736 -3364
rect 5650 -3426 5736 -3398
rect 6714 -3092 6800 -3026
rect 6714 -3126 6740 -3092
rect 6774 -3126 6800 -3092
rect 6714 -3160 6800 -3126
rect 6714 -3194 6740 -3160
rect 6774 -3194 6800 -3160
rect 6714 -3228 6800 -3194
rect 6714 -3262 6740 -3228
rect 6774 -3262 6800 -3228
rect 6714 -3296 6800 -3262
rect 6714 -3330 6740 -3296
rect 6774 -3330 6800 -3296
rect 6714 -3364 6800 -3330
rect 6714 -3398 6740 -3364
rect 6774 -3398 6800 -3364
rect 6714 -3426 6800 -3398
rect 7778 -3092 7864 -3026
rect 7778 -3126 7804 -3092
rect 7838 -3126 7864 -3092
rect 7778 -3160 7864 -3126
rect 7778 -3194 7804 -3160
rect 7838 -3194 7864 -3160
rect 7778 -3228 7864 -3194
rect 7778 -3262 7804 -3228
rect 7838 -3262 7864 -3228
rect 7778 -3296 7864 -3262
rect 7778 -3330 7804 -3296
rect 7838 -3330 7864 -3296
rect 7778 -3364 7864 -3330
rect 7778 -3398 7804 -3364
rect 7838 -3398 7864 -3364
rect 7778 -3426 7864 -3398
<< nsubdiff >>
rect 3954 470 4018 524
rect 3954 436 3958 470
rect 3992 436 4018 470
rect 3954 402 4018 436
rect 3954 368 3958 402
rect 3992 368 4018 402
rect 3954 334 4018 368
rect 3954 300 3958 334
rect 3992 300 4018 334
rect 3954 266 4018 300
rect 3954 232 3958 266
rect 3992 232 4018 266
rect 3954 198 4018 232
rect 3954 164 3958 198
rect 3992 164 4018 198
rect 3954 130 4018 164
rect 3954 96 3958 130
rect 3992 96 4018 130
rect 3954 62 4018 96
rect 3954 28 3958 62
rect 3992 28 4018 62
rect 3954 -6 4018 28
rect 3954 -40 3958 -6
rect 3992 -40 4018 -6
rect 3954 -74 4018 -40
rect 3954 -108 3958 -74
rect 3992 -108 4018 -74
rect 3954 -142 4018 -108
rect 3954 -176 3958 -142
rect 3992 -176 4018 -142
rect 3954 -210 4018 -176
rect 3954 -244 3958 -210
rect 3992 -244 4018 -210
rect 3954 -278 4018 -244
rect 3954 -312 3958 -278
rect 3992 -312 4018 -278
rect 3954 -346 4018 -312
rect 3954 -380 3958 -346
rect 3992 -380 4018 -346
rect 3954 -414 4018 -380
rect 3954 -448 3958 -414
rect 3992 -448 4018 -414
rect 3954 -476 4018 -448
rect 4996 470 5082 524
rect 4996 436 5022 470
rect 5056 436 5082 470
rect 4996 402 5082 436
rect 4996 368 5022 402
rect 5056 368 5082 402
rect 4996 334 5082 368
rect 4996 300 5022 334
rect 5056 300 5082 334
rect 4996 266 5082 300
rect 4996 232 5022 266
rect 5056 232 5082 266
rect 4996 198 5082 232
rect 4996 164 5022 198
rect 5056 164 5082 198
rect 4996 130 5082 164
rect 4996 96 5022 130
rect 5056 96 5082 130
rect 4996 62 5082 96
rect 4996 28 5022 62
rect 5056 28 5082 62
rect 4996 -6 5082 28
rect 4996 -40 5022 -6
rect 5056 -40 5082 -6
rect 4996 -74 5082 -40
rect 4996 -108 5022 -74
rect 5056 -108 5082 -74
rect 4996 -142 5082 -108
rect 4996 -176 5022 -142
rect 5056 -176 5082 -142
rect 4996 -210 5082 -176
rect 4996 -244 5022 -210
rect 5056 -244 5082 -210
rect 4996 -278 5082 -244
rect 4996 -312 5022 -278
rect 5056 -312 5082 -278
rect 4996 -346 5082 -312
rect 4996 -380 5022 -346
rect 5056 -380 5082 -346
rect 4996 -414 5082 -380
rect 4996 -448 5022 -414
rect 5056 -448 5082 -414
rect 4996 -476 5082 -448
rect 5670 470 5734 524
rect 5670 436 5674 470
rect 5708 436 5734 470
rect 5670 402 5734 436
rect 5670 368 5674 402
rect 5708 368 5734 402
rect 5670 334 5734 368
rect 5670 300 5674 334
rect 5708 300 5734 334
rect 5670 266 5734 300
rect 5670 232 5674 266
rect 5708 232 5734 266
rect 5670 198 5734 232
rect 5670 164 5674 198
rect 5708 164 5734 198
rect 5670 130 5734 164
rect 5670 96 5674 130
rect 5708 96 5734 130
rect 5670 62 5734 96
rect 5670 28 5674 62
rect 5708 28 5734 62
rect 5670 -6 5734 28
rect 5670 -40 5674 -6
rect 5708 -40 5734 -6
rect 5670 -74 5734 -40
rect 5670 -108 5674 -74
rect 5708 -108 5734 -74
rect 5670 -142 5734 -108
rect 5670 -176 5674 -142
rect 5708 -176 5734 -142
rect 5670 -210 5734 -176
rect 5670 -244 5674 -210
rect 5708 -244 5734 -210
rect 5670 -278 5734 -244
rect 5670 -312 5674 -278
rect 5708 -312 5734 -278
rect 5670 -346 5734 -312
rect 5670 -380 5674 -346
rect 5708 -380 5734 -346
rect 5670 -414 5734 -380
rect 5670 -448 5674 -414
rect 5708 -448 5734 -414
rect 5670 -476 5734 -448
rect 6712 470 6798 524
rect 6712 436 6738 470
rect 6772 436 6798 470
rect 6712 402 6798 436
rect 6712 368 6738 402
rect 6772 368 6798 402
rect 6712 334 6798 368
rect 6712 300 6738 334
rect 6772 300 6798 334
rect 6712 266 6798 300
rect 6712 232 6738 266
rect 6772 232 6798 266
rect 6712 198 6798 232
rect 6712 164 6738 198
rect 6772 164 6798 198
rect 6712 130 6798 164
rect 6712 96 6738 130
rect 6772 96 6798 130
rect 6712 62 6798 96
rect 6712 28 6738 62
rect 6772 28 6798 62
rect 6712 -6 6798 28
rect 6712 -40 6738 -6
rect 6772 -40 6798 -6
rect 6712 -74 6798 -40
rect 6712 -108 6738 -74
rect 6772 -108 6798 -74
rect 6712 -142 6798 -108
rect 6712 -176 6738 -142
rect 6772 -176 6798 -142
rect 6712 -210 6798 -176
rect 6712 -244 6738 -210
rect 6772 -244 6798 -210
rect 6712 -278 6798 -244
rect 6712 -312 6738 -278
rect 6772 -312 6798 -278
rect 6712 -346 6798 -312
rect 6712 -380 6738 -346
rect 6772 -380 6798 -346
rect 6712 -414 6798 -380
rect 6712 -448 6738 -414
rect 6772 -448 6798 -414
rect 6712 -476 6798 -448
rect 7776 470 7840 524
rect 7776 436 7802 470
rect 7836 436 7840 470
rect 7776 402 7840 436
rect 7776 368 7802 402
rect 7836 368 7840 402
rect 7776 334 7840 368
rect 7776 300 7802 334
rect 7836 300 7840 334
rect 7776 266 7840 300
rect 7776 232 7802 266
rect 7836 232 7840 266
rect 7776 198 7840 232
rect 7776 164 7802 198
rect 7836 164 7840 198
rect 7776 130 7840 164
rect 7776 96 7802 130
rect 7836 96 7840 130
rect 7776 62 7840 96
rect 7776 28 7802 62
rect 7836 28 7840 62
rect 7776 -6 7840 28
rect 7776 -40 7802 -6
rect 7836 -40 7840 -6
rect 7776 -74 7840 -40
rect 7776 -108 7802 -74
rect 7836 -108 7840 -74
rect 7776 -142 7840 -108
rect 7776 -176 7802 -142
rect 7836 -176 7840 -142
rect 7776 -210 7840 -176
rect 7776 -244 7802 -210
rect 7836 -244 7840 -210
rect 7776 -278 7840 -244
rect 7776 -312 7802 -278
rect 7836 -312 7840 -278
rect 7776 -346 7840 -312
rect 7776 -380 7802 -346
rect 7836 -380 7840 -346
rect 7776 -414 7840 -380
rect 7776 -448 7802 -414
rect 7836 -448 7840 -414
rect 7776 -476 7840 -448
rect 3954 -1438 4018 -1384
rect 3954 -1472 3958 -1438
rect 3992 -1472 4018 -1438
rect 3954 -1506 4018 -1472
rect 3954 -1540 3958 -1506
rect 3992 -1540 4018 -1506
rect 3954 -1574 4018 -1540
rect 3954 -1608 3958 -1574
rect 3992 -1608 4018 -1574
rect 3954 -1642 4018 -1608
rect 3954 -1676 3958 -1642
rect 3992 -1676 4018 -1642
rect 3954 -1710 4018 -1676
rect 3954 -1744 3958 -1710
rect 3992 -1744 4018 -1710
rect 3954 -1778 4018 -1744
rect 3954 -1812 3958 -1778
rect 3992 -1812 4018 -1778
rect 3954 -1846 4018 -1812
rect 3954 -1880 3958 -1846
rect 3992 -1880 4018 -1846
rect 3954 -1914 4018 -1880
rect 3954 -1948 3958 -1914
rect 3992 -1948 4018 -1914
rect 3954 -1982 4018 -1948
rect 3954 -2016 3958 -1982
rect 3992 -2016 4018 -1982
rect 3954 -2050 4018 -2016
rect 3954 -2084 3958 -2050
rect 3992 -2084 4018 -2050
rect 3954 -2118 4018 -2084
rect 3954 -2152 3958 -2118
rect 3992 -2152 4018 -2118
rect 3954 -2186 4018 -2152
rect 3954 -2220 3958 -2186
rect 3992 -2220 4018 -2186
rect 3954 -2254 4018 -2220
rect 3954 -2288 3958 -2254
rect 3992 -2288 4018 -2254
rect 3954 -2322 4018 -2288
rect 3954 -2356 3958 -2322
rect 3992 -2356 4018 -2322
rect 3954 -2384 4018 -2356
rect 4996 -1438 5082 -1384
rect 4996 -1472 5022 -1438
rect 5056 -1472 5082 -1438
rect 4996 -1506 5082 -1472
rect 4996 -1540 5022 -1506
rect 5056 -1540 5082 -1506
rect 4996 -1574 5082 -1540
rect 4996 -1608 5022 -1574
rect 5056 -1608 5082 -1574
rect 4996 -1642 5082 -1608
rect 4996 -1676 5022 -1642
rect 5056 -1676 5082 -1642
rect 4996 -1710 5082 -1676
rect 4996 -1744 5022 -1710
rect 5056 -1744 5082 -1710
rect 4996 -1778 5082 -1744
rect 4996 -1812 5022 -1778
rect 5056 -1812 5082 -1778
rect 4996 -1846 5082 -1812
rect 4996 -1880 5022 -1846
rect 5056 -1880 5082 -1846
rect 4996 -1914 5082 -1880
rect 4996 -1948 5022 -1914
rect 5056 -1948 5082 -1914
rect 4996 -1982 5082 -1948
rect 4996 -2016 5022 -1982
rect 5056 -2016 5082 -1982
rect 4996 -2050 5082 -2016
rect 4996 -2084 5022 -2050
rect 5056 -2084 5082 -2050
rect 4996 -2118 5082 -2084
rect 4996 -2152 5022 -2118
rect 5056 -2152 5082 -2118
rect 4996 -2186 5082 -2152
rect 4996 -2220 5022 -2186
rect 5056 -2220 5082 -2186
rect 4996 -2254 5082 -2220
rect 4996 -2288 5022 -2254
rect 5056 -2288 5082 -2254
rect 4996 -2322 5082 -2288
rect 4996 -2356 5022 -2322
rect 5056 -2356 5082 -2322
rect 4996 -2384 5082 -2356
rect 5672 -1438 5736 -1384
rect 5672 -1472 5676 -1438
rect 5710 -1472 5736 -1438
rect 5672 -1506 5736 -1472
rect 5672 -1540 5676 -1506
rect 5710 -1540 5736 -1506
rect 5672 -1574 5736 -1540
rect 5672 -1608 5676 -1574
rect 5710 -1608 5736 -1574
rect 5672 -1642 5736 -1608
rect 5672 -1676 5676 -1642
rect 5710 -1676 5736 -1642
rect 5672 -1710 5736 -1676
rect 5672 -1744 5676 -1710
rect 5710 -1744 5736 -1710
rect 5672 -1778 5736 -1744
rect 5672 -1812 5676 -1778
rect 5710 -1812 5736 -1778
rect 5672 -1846 5736 -1812
rect 5672 -1880 5676 -1846
rect 5710 -1880 5736 -1846
rect 5672 -1914 5736 -1880
rect 5672 -1948 5676 -1914
rect 5710 -1948 5736 -1914
rect 5672 -1982 5736 -1948
rect 5672 -2016 5676 -1982
rect 5710 -2016 5736 -1982
rect 5672 -2050 5736 -2016
rect 5672 -2084 5676 -2050
rect 5710 -2084 5736 -2050
rect 5672 -2118 5736 -2084
rect 5672 -2152 5676 -2118
rect 5710 -2152 5736 -2118
rect 5672 -2186 5736 -2152
rect 5672 -2220 5676 -2186
rect 5710 -2220 5736 -2186
rect 5672 -2254 5736 -2220
rect 5672 -2288 5676 -2254
rect 5710 -2288 5736 -2254
rect 5672 -2322 5736 -2288
rect 5672 -2356 5676 -2322
rect 5710 -2356 5736 -2322
rect 5672 -2384 5736 -2356
rect 6714 -1438 6800 -1384
rect 6714 -1472 6740 -1438
rect 6774 -1472 6800 -1438
rect 6714 -1506 6800 -1472
rect 6714 -1540 6740 -1506
rect 6774 -1540 6800 -1506
rect 6714 -1574 6800 -1540
rect 6714 -1608 6740 -1574
rect 6774 -1608 6800 -1574
rect 6714 -1642 6800 -1608
rect 6714 -1676 6740 -1642
rect 6774 -1676 6800 -1642
rect 6714 -1710 6800 -1676
rect 6714 -1744 6740 -1710
rect 6774 -1744 6800 -1710
rect 6714 -1778 6800 -1744
rect 6714 -1812 6740 -1778
rect 6774 -1812 6800 -1778
rect 6714 -1846 6800 -1812
rect 6714 -1880 6740 -1846
rect 6774 -1880 6800 -1846
rect 6714 -1914 6800 -1880
rect 6714 -1948 6740 -1914
rect 6774 -1948 6800 -1914
rect 6714 -1982 6800 -1948
rect 6714 -2016 6740 -1982
rect 6774 -2016 6800 -1982
rect 6714 -2050 6800 -2016
rect 6714 -2084 6740 -2050
rect 6774 -2084 6800 -2050
rect 6714 -2118 6800 -2084
rect 6714 -2152 6740 -2118
rect 6774 -2152 6800 -2118
rect 6714 -2186 6800 -2152
rect 6714 -2220 6740 -2186
rect 6774 -2220 6800 -2186
rect 6714 -2254 6800 -2220
rect 6714 -2288 6740 -2254
rect 6774 -2288 6800 -2254
rect 6714 -2322 6800 -2288
rect 6714 -2356 6740 -2322
rect 6774 -2356 6800 -2322
rect 6714 -2384 6800 -2356
rect 7778 -1438 7842 -1384
rect 7778 -1472 7804 -1438
rect 7838 -1472 7842 -1438
rect 7778 -1506 7842 -1472
rect 7778 -1540 7804 -1506
rect 7838 -1540 7842 -1506
rect 7778 -1574 7842 -1540
rect 7778 -1608 7804 -1574
rect 7838 -1608 7842 -1574
rect 7778 -1642 7842 -1608
rect 7778 -1676 7804 -1642
rect 7838 -1676 7842 -1642
rect 7778 -1710 7842 -1676
rect 7778 -1744 7804 -1710
rect 7838 -1744 7842 -1710
rect 7778 -1778 7842 -1744
rect 7778 -1812 7804 -1778
rect 7838 -1812 7842 -1778
rect 7778 -1846 7842 -1812
rect 7778 -1880 7804 -1846
rect 7838 -1880 7842 -1846
rect 7778 -1914 7842 -1880
rect 7778 -1948 7804 -1914
rect 7838 -1948 7842 -1914
rect 7778 -1982 7842 -1948
rect 7778 -2016 7804 -1982
rect 7838 -2016 7842 -1982
rect 7778 -2050 7842 -2016
rect 7778 -2084 7804 -2050
rect 7838 -2084 7842 -2050
rect 7778 -2118 7842 -2084
rect 7778 -2152 7804 -2118
rect 7838 -2152 7842 -2118
rect 7778 -2186 7842 -2152
rect 7778 -2220 7804 -2186
rect 7838 -2220 7842 -2186
rect 7778 -2254 7842 -2220
rect 7778 -2288 7804 -2254
rect 7838 -2288 7842 -2254
rect 7778 -2322 7842 -2288
rect 7778 -2356 7804 -2322
rect 7838 -2356 7842 -2322
rect 7778 -2384 7842 -2356
<< psubdiffcont >>
rect 3548 -3126 3582 -3092
rect 3548 -3194 3582 -3160
rect 3548 -3262 3582 -3228
rect 3548 -3330 3582 -3296
rect 3548 -3398 3582 -3364
rect 4612 -3126 4646 -3092
rect 4612 -3194 4646 -3160
rect 4612 -3262 4646 -3228
rect 4612 -3330 4646 -3296
rect 4612 -3398 4646 -3364
rect 5676 -3126 5710 -3092
rect 5676 -3194 5710 -3160
rect 5676 -3262 5710 -3228
rect 5676 -3330 5710 -3296
rect 5676 -3398 5710 -3364
rect 6740 -3126 6774 -3092
rect 6740 -3194 6774 -3160
rect 6740 -3262 6774 -3228
rect 6740 -3330 6774 -3296
rect 6740 -3398 6774 -3364
rect 7804 -3126 7838 -3092
rect 7804 -3194 7838 -3160
rect 7804 -3262 7838 -3228
rect 7804 -3330 7838 -3296
rect 7804 -3398 7838 -3364
<< nsubdiffcont >>
rect 3958 436 3992 470
rect 3958 368 3992 402
rect 3958 300 3992 334
rect 3958 232 3992 266
rect 3958 164 3992 198
rect 3958 96 3992 130
rect 3958 28 3992 62
rect 3958 -40 3992 -6
rect 3958 -108 3992 -74
rect 3958 -176 3992 -142
rect 3958 -244 3992 -210
rect 3958 -312 3992 -278
rect 3958 -380 3992 -346
rect 3958 -448 3992 -414
rect 5022 436 5056 470
rect 5022 368 5056 402
rect 5022 300 5056 334
rect 5022 232 5056 266
rect 5022 164 5056 198
rect 5022 96 5056 130
rect 5022 28 5056 62
rect 5022 -40 5056 -6
rect 5022 -108 5056 -74
rect 5022 -176 5056 -142
rect 5022 -244 5056 -210
rect 5022 -312 5056 -278
rect 5022 -380 5056 -346
rect 5022 -448 5056 -414
rect 5674 436 5708 470
rect 5674 368 5708 402
rect 5674 300 5708 334
rect 5674 232 5708 266
rect 5674 164 5708 198
rect 5674 96 5708 130
rect 5674 28 5708 62
rect 5674 -40 5708 -6
rect 5674 -108 5708 -74
rect 5674 -176 5708 -142
rect 5674 -244 5708 -210
rect 5674 -312 5708 -278
rect 5674 -380 5708 -346
rect 5674 -448 5708 -414
rect 6738 436 6772 470
rect 6738 368 6772 402
rect 6738 300 6772 334
rect 6738 232 6772 266
rect 6738 164 6772 198
rect 6738 96 6772 130
rect 6738 28 6772 62
rect 6738 -40 6772 -6
rect 6738 -108 6772 -74
rect 6738 -176 6772 -142
rect 6738 -244 6772 -210
rect 6738 -312 6772 -278
rect 6738 -380 6772 -346
rect 6738 -448 6772 -414
rect 7802 436 7836 470
rect 7802 368 7836 402
rect 7802 300 7836 334
rect 7802 232 7836 266
rect 7802 164 7836 198
rect 7802 96 7836 130
rect 7802 28 7836 62
rect 7802 -40 7836 -6
rect 7802 -108 7836 -74
rect 7802 -176 7836 -142
rect 7802 -244 7836 -210
rect 7802 -312 7836 -278
rect 7802 -380 7836 -346
rect 7802 -448 7836 -414
rect 3958 -1472 3992 -1438
rect 3958 -1540 3992 -1506
rect 3958 -1608 3992 -1574
rect 3958 -1676 3992 -1642
rect 3958 -1744 3992 -1710
rect 3958 -1812 3992 -1778
rect 3958 -1880 3992 -1846
rect 3958 -1948 3992 -1914
rect 3958 -2016 3992 -1982
rect 3958 -2084 3992 -2050
rect 3958 -2152 3992 -2118
rect 3958 -2220 3992 -2186
rect 3958 -2288 3992 -2254
rect 3958 -2356 3992 -2322
rect 5022 -1472 5056 -1438
rect 5022 -1540 5056 -1506
rect 5022 -1608 5056 -1574
rect 5022 -1676 5056 -1642
rect 5022 -1744 5056 -1710
rect 5022 -1812 5056 -1778
rect 5022 -1880 5056 -1846
rect 5022 -1948 5056 -1914
rect 5022 -2016 5056 -1982
rect 5022 -2084 5056 -2050
rect 5022 -2152 5056 -2118
rect 5022 -2220 5056 -2186
rect 5022 -2288 5056 -2254
rect 5022 -2356 5056 -2322
rect 5676 -1472 5710 -1438
rect 5676 -1540 5710 -1506
rect 5676 -1608 5710 -1574
rect 5676 -1676 5710 -1642
rect 5676 -1744 5710 -1710
rect 5676 -1812 5710 -1778
rect 5676 -1880 5710 -1846
rect 5676 -1948 5710 -1914
rect 5676 -2016 5710 -1982
rect 5676 -2084 5710 -2050
rect 5676 -2152 5710 -2118
rect 5676 -2220 5710 -2186
rect 5676 -2288 5710 -2254
rect 5676 -2356 5710 -2322
rect 6740 -1472 6774 -1438
rect 6740 -1540 6774 -1506
rect 6740 -1608 6774 -1574
rect 6740 -1676 6774 -1642
rect 6740 -1744 6774 -1710
rect 6740 -1812 6774 -1778
rect 6740 -1880 6774 -1846
rect 6740 -1948 6774 -1914
rect 6740 -2016 6774 -1982
rect 6740 -2084 6774 -2050
rect 6740 -2152 6774 -2118
rect 6740 -2220 6774 -2186
rect 6740 -2288 6774 -2254
rect 6740 -2356 6774 -2322
rect 7804 -1472 7838 -1438
rect 7804 -1540 7838 -1506
rect 7804 -1608 7838 -1574
rect 7804 -1676 7838 -1642
rect 7804 -1744 7838 -1710
rect 7804 -1812 7838 -1778
rect 7804 -1880 7838 -1846
rect 7804 -1948 7838 -1914
rect 7804 -2016 7838 -1982
rect 7804 -2084 7838 -2050
rect 7804 -2152 7838 -2118
rect 7804 -2220 7838 -2186
rect 7804 -2288 7838 -2254
rect 7804 -2356 7838 -2322
<< locali >>
rect 3958 512 3992 528
rect 3958 -480 3992 -464
rect 5022 512 5056 528
rect 5022 -480 5056 -464
rect 5674 512 5708 528
rect 6738 512 6772 528
rect 6206 22 6240 30
rect 5674 -480 5708 -464
rect 6738 -480 6772 -464
rect 7802 512 7836 528
rect 7802 -480 7836 -464
rect 3958 -1396 3992 -1380
rect 3958 -2388 3992 -2372
rect 5022 -1396 5056 -1380
rect 5022 -2388 5056 -2372
rect 5676 -1396 5710 -1380
rect 6208 -1402 6242 -1394
rect 6740 -1396 6774 -1380
rect 5676 -2388 5710 -2372
rect 6740 -2388 6774 -2372
rect 7804 -1396 7838 -1380
rect 7804 -2388 7838 -2372
rect 3548 -3038 3582 -3022
rect 3548 -3430 3582 -3414
rect 4612 -3038 4646 -3022
rect 4612 -3430 4646 -3414
rect 5676 -3038 5710 -3022
rect 5676 -3430 5710 -3414
rect 6740 -3038 6774 -3022
rect 6740 -3430 6774 -3414
rect 7804 -3038 7838 -3022
rect 7804 -3430 7838 -3414
<< viali >>
rect 3958 470 3992 512
rect 3958 436 3992 470
rect 3958 402 3992 436
rect 3958 368 3992 402
rect 3958 334 3992 368
rect 3958 300 3992 334
rect 3958 266 3992 300
rect 3958 232 3992 266
rect 3958 198 3992 232
rect 3958 164 3992 198
rect 3958 130 3992 164
rect 3958 96 3992 130
rect 3958 62 3992 96
rect 3958 28 3992 62
rect 3958 -6 3992 28
rect 3958 -40 3992 -6
rect 3958 -74 3992 -40
rect 3958 -108 3992 -74
rect 3958 -142 3992 -108
rect 3958 -176 3992 -142
rect 3958 -210 3992 -176
rect 3958 -244 3992 -210
rect 3958 -278 3992 -244
rect 3958 -312 3992 -278
rect 3958 -346 3992 -312
rect 3958 -380 3992 -346
rect 3958 -414 3992 -380
rect 3958 -448 3992 -414
rect 3958 -464 3992 -448
rect 5022 470 5056 512
rect 5022 436 5056 470
rect 5022 402 5056 436
rect 5022 368 5056 402
rect 5022 334 5056 368
rect 5022 300 5056 334
rect 5022 266 5056 300
rect 5022 232 5056 266
rect 5022 198 5056 232
rect 5022 164 5056 198
rect 5022 130 5056 164
rect 5022 96 5056 130
rect 5022 62 5056 96
rect 5022 28 5056 62
rect 5022 -6 5056 28
rect 5022 -40 5056 -6
rect 5022 -74 5056 -40
rect 5022 -108 5056 -74
rect 5022 -142 5056 -108
rect 5022 -176 5056 -142
rect 5022 -210 5056 -176
rect 5022 -244 5056 -210
rect 5022 -278 5056 -244
rect 5022 -312 5056 -278
rect 5022 -346 5056 -312
rect 5022 -380 5056 -346
rect 5022 -414 5056 -380
rect 5022 -448 5056 -414
rect 5022 -464 5056 -448
rect 5674 470 5708 512
rect 5674 436 5708 470
rect 5674 402 5708 436
rect 5674 368 5708 402
rect 5674 334 5708 368
rect 5674 300 5708 334
rect 5674 266 5708 300
rect 5674 232 5708 266
rect 5674 198 5708 232
rect 5674 164 5708 198
rect 5674 130 5708 164
rect 5674 96 5708 130
rect 5674 62 5708 96
rect 5674 28 5708 62
rect 6738 470 6772 512
rect 6738 436 6772 470
rect 6738 402 6772 436
rect 6738 368 6772 402
rect 6738 334 6772 368
rect 6738 300 6772 334
rect 6738 266 6772 300
rect 6738 232 6772 266
rect 6738 198 6772 232
rect 6738 164 6772 198
rect 6738 130 6772 164
rect 6738 96 6772 130
rect 6738 62 6772 96
rect 5674 -6 5708 28
rect 6738 28 6772 62
rect 5674 -40 5708 -6
rect 5674 -74 5708 -40
rect 5674 -108 5708 -74
rect 5674 -142 5708 -108
rect 5674 -176 5708 -142
rect 5674 -210 5708 -176
rect 5674 -244 5708 -210
rect 5674 -278 5708 -244
rect 5674 -312 5708 -278
rect 5674 -346 5708 -312
rect 5674 -380 5708 -346
rect 5674 -414 5708 -380
rect 5674 -448 5708 -414
rect 5674 -464 5708 -448
rect 6738 -6 6772 28
rect 6738 -40 6772 -6
rect 6738 -74 6772 -40
rect 6738 -108 6772 -74
rect 6738 -142 6772 -108
rect 6738 -176 6772 -142
rect 6738 -210 6772 -176
rect 6738 -244 6772 -210
rect 6738 -278 6772 -244
rect 6738 -312 6772 -278
rect 6738 -346 6772 -312
rect 6738 -380 6772 -346
rect 6738 -414 6772 -380
rect 6738 -448 6772 -414
rect 6738 -464 6772 -448
rect 7802 470 7836 512
rect 7802 436 7836 470
rect 7802 402 7836 436
rect 7802 368 7836 402
rect 7802 334 7836 368
rect 7802 300 7836 334
rect 7802 266 7836 300
rect 7802 232 7836 266
rect 7802 198 7836 232
rect 7802 164 7836 198
rect 7802 130 7836 164
rect 7802 96 7836 130
rect 7802 62 7836 96
rect 7802 28 7836 62
rect 7802 -6 7836 28
rect 7802 -40 7836 -6
rect 7802 -74 7836 -40
rect 7802 -108 7836 -74
rect 7802 -142 7836 -108
rect 7802 -176 7836 -142
rect 7802 -210 7836 -176
rect 7802 -244 7836 -210
rect 7802 -278 7836 -244
rect 7802 -312 7836 -278
rect 7802 -346 7836 -312
rect 7802 -380 7836 -346
rect 7802 -414 7836 -380
rect 7802 -448 7836 -414
rect 7802 -464 7836 -448
rect 3958 -1438 3992 -1396
rect 3958 -1472 3992 -1438
rect 3958 -1506 3992 -1472
rect 3958 -1540 3992 -1506
rect 3958 -1574 3992 -1540
rect 3958 -1608 3992 -1574
rect 3958 -1642 3992 -1608
rect 3958 -1676 3992 -1642
rect 3958 -1710 3992 -1676
rect 3958 -1744 3992 -1710
rect 3958 -1778 3992 -1744
rect 3958 -1812 3992 -1778
rect 3958 -1846 3992 -1812
rect 3958 -1880 3992 -1846
rect 3958 -1914 3992 -1880
rect 3958 -1948 3992 -1914
rect 3958 -1982 3992 -1948
rect 3958 -2016 3992 -1982
rect 3958 -2050 3992 -2016
rect 3958 -2084 3992 -2050
rect 3958 -2118 3992 -2084
rect 3958 -2152 3992 -2118
rect 3958 -2186 3992 -2152
rect 3958 -2220 3992 -2186
rect 3958 -2254 3992 -2220
rect 3958 -2288 3992 -2254
rect 3958 -2322 3992 -2288
rect 3958 -2356 3992 -2322
rect 3958 -2372 3992 -2356
rect 5022 -1438 5056 -1396
rect 5022 -1472 5056 -1438
rect 5022 -1506 5056 -1472
rect 5022 -1540 5056 -1506
rect 5022 -1574 5056 -1540
rect 5022 -1608 5056 -1574
rect 5022 -1642 5056 -1608
rect 5022 -1676 5056 -1642
rect 5022 -1710 5056 -1676
rect 5022 -1744 5056 -1710
rect 5022 -1778 5056 -1744
rect 5022 -1812 5056 -1778
rect 5022 -1846 5056 -1812
rect 5022 -1880 5056 -1846
rect 5022 -1914 5056 -1880
rect 5022 -1948 5056 -1914
rect 5022 -1982 5056 -1948
rect 5022 -2016 5056 -1982
rect 5022 -2050 5056 -2016
rect 5022 -2084 5056 -2050
rect 5022 -2118 5056 -2084
rect 5022 -2152 5056 -2118
rect 5022 -2186 5056 -2152
rect 5022 -2220 5056 -2186
rect 5022 -2254 5056 -2220
rect 5022 -2288 5056 -2254
rect 5022 -2322 5056 -2288
rect 5022 -2356 5056 -2322
rect 5022 -2372 5056 -2356
rect 5676 -1438 5710 -1396
rect 5676 -1472 5710 -1438
rect 5676 -1506 5710 -1472
rect 5676 -1540 5710 -1506
rect 5676 -1574 5710 -1540
rect 5676 -1608 5710 -1574
rect 5676 -1642 5710 -1608
rect 5676 -1676 5710 -1642
rect 5676 -1710 5710 -1676
rect 5676 -1744 5710 -1710
rect 5676 -1778 5710 -1744
rect 5676 -1812 5710 -1778
rect 5676 -1846 5710 -1812
rect 5676 -1880 5710 -1846
rect 5676 -1914 5710 -1880
rect 5676 -1948 5710 -1914
rect 5676 -1982 5710 -1948
rect 5676 -2016 5710 -1982
rect 5676 -2050 5710 -2016
rect 5676 -2084 5710 -2050
rect 5676 -2118 5710 -2084
rect 5676 -2152 5710 -2118
rect 5676 -2186 5710 -2152
rect 5676 -2220 5710 -2186
rect 5676 -2254 5710 -2220
rect 5676 -2288 5710 -2254
rect 5676 -2322 5710 -2288
rect 5676 -2356 5710 -2322
rect 5676 -2372 5710 -2356
rect 6740 -1438 6774 -1396
rect 6740 -1472 6774 -1438
rect 6740 -1506 6774 -1472
rect 6740 -1540 6774 -1506
rect 6740 -1574 6774 -1540
rect 6740 -1608 6774 -1574
rect 6740 -1642 6774 -1608
rect 6740 -1676 6774 -1642
rect 6740 -1710 6774 -1676
rect 6740 -1744 6774 -1710
rect 6740 -1778 6774 -1744
rect 6740 -1812 6774 -1778
rect 6740 -1846 6774 -1812
rect 6740 -1880 6774 -1846
rect 6740 -1914 6774 -1880
rect 6740 -1948 6774 -1914
rect 6740 -1982 6774 -1948
rect 6740 -2016 6774 -1982
rect 6740 -2050 6774 -2016
rect 6740 -2084 6774 -2050
rect 6740 -2118 6774 -2084
rect 6740 -2152 6774 -2118
rect 6740 -2186 6774 -2152
rect 6740 -2220 6774 -2186
rect 6740 -2254 6774 -2220
rect 6740 -2288 6774 -2254
rect 6740 -2322 6774 -2288
rect 6740 -2356 6774 -2322
rect 6740 -2372 6774 -2356
rect 7804 -1438 7838 -1396
rect 7804 -1472 7838 -1438
rect 7804 -1506 7838 -1472
rect 7804 -1540 7838 -1506
rect 7804 -1574 7838 -1540
rect 7804 -1608 7838 -1574
rect 7804 -1642 7838 -1608
rect 7804 -1676 7838 -1642
rect 7804 -1710 7838 -1676
rect 7804 -1744 7838 -1710
rect 7804 -1778 7838 -1744
rect 7804 -1812 7838 -1778
rect 7804 -1846 7838 -1812
rect 7804 -1880 7838 -1846
rect 7804 -1914 7838 -1880
rect 7804 -1948 7838 -1914
rect 7804 -1982 7838 -1948
rect 7804 -2016 7838 -1982
rect 7804 -2050 7838 -2016
rect 7804 -2084 7838 -2050
rect 7804 -2118 7838 -2084
rect 7804 -2152 7838 -2118
rect 7804 -2186 7838 -2152
rect 7804 -2220 7838 -2186
rect 7804 -2254 7838 -2220
rect 7804 -2288 7838 -2254
rect 7804 -2322 7838 -2288
rect 7804 -2356 7838 -2322
rect 7804 -2372 7838 -2356
rect 3548 -3092 3582 -3038
rect 3548 -3126 3582 -3092
rect 3548 -3160 3582 -3126
rect 3548 -3194 3582 -3160
rect 3548 -3228 3582 -3194
rect 3548 -3262 3582 -3228
rect 3548 -3296 3582 -3262
rect 3548 -3330 3582 -3296
rect 3548 -3364 3582 -3330
rect 3548 -3398 3582 -3364
rect 3548 -3414 3582 -3398
rect 4612 -3092 4646 -3038
rect 4612 -3126 4646 -3092
rect 4612 -3160 4646 -3126
rect 4612 -3194 4646 -3160
rect 4612 -3228 4646 -3194
rect 4612 -3262 4646 -3228
rect 4612 -3296 4646 -3262
rect 4612 -3330 4646 -3296
rect 4612 -3364 4646 -3330
rect 4612 -3398 4646 -3364
rect 4612 -3414 4646 -3398
rect 5676 -3092 5710 -3038
rect 5676 -3126 5710 -3092
rect 5676 -3160 5710 -3126
rect 5676 -3194 5710 -3160
rect 5676 -3228 5710 -3194
rect 5676 -3262 5710 -3228
rect 5676 -3296 5710 -3262
rect 5676 -3330 5710 -3296
rect 5676 -3364 5710 -3330
rect 5676 -3398 5710 -3364
rect 5676 -3414 5710 -3398
rect 6740 -3092 6774 -3038
rect 6740 -3126 6774 -3092
rect 6740 -3160 6774 -3126
rect 6740 -3194 6774 -3160
rect 6740 -3228 6774 -3194
rect 6740 -3262 6774 -3228
rect 6740 -3296 6774 -3262
rect 6740 -3330 6774 -3296
rect 6740 -3364 6774 -3330
rect 6740 -3398 6774 -3364
rect 6740 -3414 6774 -3398
rect 7804 -3092 7838 -3038
rect 7804 -3126 7838 -3092
rect 7804 -3160 7838 -3126
rect 7804 -3194 7838 -3160
rect 7804 -3228 7838 -3194
rect 7804 -3262 7838 -3228
rect 7804 -3296 7838 -3262
rect 7804 -3330 7838 -3296
rect 7804 -3364 7838 -3330
rect 7804 -3398 7838 -3364
rect 7804 -3414 7838 -3398
<< metal1 >>
rect 3946 3226 4050 3232
rect 3336 -594 3588 542
rect 3946 512 4050 2776
rect 4988 3226 5092 3232
rect 4988 524 5092 2776
rect 5636 3226 5740 3232
rect 5636 2770 5740 2776
rect 6704 3226 6808 3232
rect 6704 2770 6808 2776
rect 7798 3226 7902 3232
rect 5566 692 5624 698
rect 3946 -464 3958 512
rect 3992 -464 4050 512
rect 3336 -706 3342 -594
rect 3582 -706 3588 -594
rect 3336 -752 3588 -706
rect 3740 -566 3746 -514
rect 3838 -566 3844 -514
rect 3336 -1014 3588 -968
rect 3336 -1126 3342 -1014
rect 3582 -1126 3588 -1014
rect 3336 -2262 3588 -1126
rect 3740 -2946 3844 -566
rect 3946 -1396 4050 -464
rect 4478 -514 4536 524
rect 4942 512 5136 524
rect 5566 520 5624 592
rect 4942 -464 5022 512
rect 5056 -464 5136 512
rect 5534 514 5624 520
rect 5588 24 5624 514
rect 5534 18 5624 24
rect 4942 -476 5136 -464
rect 4088 -566 4094 -514
rect 4920 -566 4926 -514
rect 4546 -1294 4926 -566
rect 4088 -1346 4094 -1294
rect 4462 -1346 4468 -1294
rect 4546 -1346 4552 -1294
rect 4920 -1346 4926 -1294
rect 4988 -1384 5092 -476
rect 5152 -566 5158 -514
rect 5526 -566 5532 -514
rect 5152 -1346 5158 -1294
rect 5526 -1346 5532 -1294
rect 3946 -2372 3958 -1396
rect 3992 -2372 4050 -1396
rect 3946 -2384 4050 -2372
rect 4478 -2672 4536 -1384
rect 4942 -1396 5136 -1384
rect 4942 -2372 5022 -1396
rect 5056 -2372 5136 -1396
rect 5566 -1876 5624 18
rect 4942 -2384 5136 -2372
rect 5536 -1882 5624 -1876
rect 5588 -2372 5624 -1882
rect 5536 -2378 5624 -2372
rect 5566 -2532 5624 -2378
rect 5658 512 5714 2770
rect 6644 692 6702 698
rect 5658 -464 5674 512
rect 5708 -464 5714 512
rect 5748 512 5802 518
rect 6644 512 6702 592
rect 5748 16 5802 22
rect 6198 24 6250 30
rect 5658 -1384 5714 -464
rect 6698 406 6702 512
rect 6732 512 6778 2770
rect 7708 692 7766 698
rect 6644 16 6698 22
rect 6198 -470 6206 -464
rect 6200 -476 6206 -470
rect 6240 -470 6250 -464
rect 6732 -464 6738 512
rect 6772 -464 6778 512
rect 6812 512 6866 518
rect 7264 30 7270 34
rect 6812 16 6866 22
rect 7262 24 7270 30
rect 7304 30 7310 34
rect 7304 24 7314 30
rect 6240 -476 6246 -470
rect 6732 -476 6778 -464
rect 7262 -470 7314 -464
rect 7264 -476 7310 -470
rect 7708 -476 7766 592
rect 7798 524 7902 2776
rect 9420 1146 9672 2130
rect 9420 1030 9426 1146
rect 9666 1030 9672 1146
rect 9420 836 9672 1030
rect 7796 512 7902 524
rect 7796 -464 7802 512
rect 7836 -464 7902 512
rect 7796 -476 7902 -464
rect 5804 -566 5810 -514
rect 6178 -566 6184 -514
rect 6262 -566 6268 -514
rect 6636 -566 6642 -514
rect 5804 -594 6184 -566
rect 5804 -706 5810 -594
rect 6178 -706 6184 -594
rect 5806 -1126 5812 -1014
rect 6180 -1126 6186 -1014
rect 5806 -1294 6182 -1126
rect 5806 -1346 5812 -1294
rect 6180 -1346 6186 -1294
rect 6264 -1346 6270 -1294
rect 6638 -1346 6644 -1294
rect 6734 -1350 6778 -476
rect 6868 -566 6874 -514
rect 7242 -566 7332 -514
rect 7700 -566 7706 -514
rect 7326 -594 7706 -566
rect 6868 -706 6874 -594
rect 7242 -706 7248 -594
rect 7326 -706 7332 -594
rect 7700 -706 7706 -594
rect 6870 -1154 7248 -706
rect 7328 -1014 7706 -706
rect 7328 -1126 7334 -1014
rect 7702 -1126 7708 -1014
rect 6870 -1266 6876 -1154
rect 7244 -1266 7250 -1154
rect 6870 -1294 7250 -1266
rect 6870 -1346 6876 -1294
rect 7244 -1346 7250 -1294
rect 7328 -1346 7334 -1294
rect 7702 -1346 7708 -1294
rect 5658 -1396 5716 -1384
rect 5658 -2372 5676 -1396
rect 5710 -2372 5716 -1396
rect 6200 -1400 6252 -1394
rect 5658 -2384 5716 -2372
rect 5750 -1882 5802 -1876
rect 6734 -1396 6780 -1350
rect 6200 -1894 6208 -1888
rect 6202 -1900 6208 -1894
rect 6242 -1894 6252 -1888
rect 6646 -1882 6700 -1876
rect 6242 -1900 6248 -1894
rect 5750 -2378 5802 -2372
rect 6700 -2372 6704 -2368
rect 5566 -2638 5624 -2632
rect 6646 -2532 6704 -2372
rect 6734 -2372 6740 -1396
rect 6774 -2372 6780 -1396
rect 7264 -1394 7316 -1388
rect 6734 -2384 6780 -2372
rect 6814 -1882 6868 -1876
rect 6814 -2378 6868 -2372
rect 7260 -1882 7264 -1870
rect 7316 -1882 7318 -1870
rect 6646 -2638 6704 -2632
rect 4478 -2778 4536 -2772
rect 5132 -2812 5190 -2806
rect 5132 -2946 5190 -2912
rect 7260 -2812 7318 -1882
rect 7708 -2532 7766 -1384
rect 7798 -1396 7902 -476
rect 7798 -2372 7804 -1396
rect 7838 -2372 7902 -1396
rect 7798 -2384 7902 -2372
rect 7708 -2638 7766 -2632
rect 7260 -2918 7318 -2912
rect 8324 -2672 8382 -2666
rect 3678 -2998 3684 -2946
rect 4510 -2998 4516 -2946
rect 4742 -2998 4748 -2946
rect 5574 -2998 5580 -2946
rect 5806 -2998 5812 -2946
rect 6180 -2998 6186 -2946
rect 6264 -2998 6270 -2946
rect 6638 -2998 6644 -2946
rect 3542 -3038 3662 -3026
rect 3542 -3414 3548 -3038
rect 3582 -3414 3662 -3038
rect 3542 -4634 3662 -3414
rect 4068 -3426 4126 -2998
rect 4532 -3038 4726 -3026
rect 4532 -3414 4612 -3038
rect 4646 -3414 4726 -3038
rect 3542 -5096 3662 -5090
rect 4532 -4634 4726 -3414
rect 5132 -3426 5190 -2998
rect 5596 -3038 5790 -3026
rect 5596 -3414 5676 -3038
rect 5710 -3414 5790 -3038
rect 4532 -5096 4726 -5090
rect 5596 -4634 5790 -3414
rect 6200 -3038 6252 -3032
rect 6200 -3420 6252 -3414
rect 6660 -3038 6854 -3026
rect 6660 -3414 6740 -3038
rect 6774 -3414 6854 -3038
rect 5596 -5096 5790 -5090
rect 6660 -3426 6854 -3414
rect 7264 -3038 7316 -3032
rect 7264 -3420 7316 -3414
rect 7724 -3038 7918 -3026
rect 7724 -3414 7804 -3038
rect 7838 -3414 7918 -3038
rect 7724 -3426 7918 -3414
rect 8324 -3038 8382 -2772
rect 8324 -3414 8328 -3038
rect 8380 -3414 8382 -3038
rect 8324 -3426 8382 -3414
rect 6660 -4634 6836 -3426
rect 6870 -3506 6876 -3454
rect 7244 -3506 7250 -3454
rect 7328 -3506 7334 -3454
rect 7702 -3506 7708 -3454
rect 6660 -5096 6836 -5090
rect 7746 -4634 7896 -3426
rect 7934 -3506 7940 -3454
rect 8308 -3506 8314 -3454
rect 7746 -5096 7896 -5090
<< via1 >>
rect 3946 2776 4050 3226
rect 4988 2776 5092 3226
rect 5636 2776 5740 3226
rect 6704 2776 6808 3226
rect 7798 2776 7902 3226
rect 5566 592 5624 692
rect 3342 -706 3582 -594
rect 3746 -566 3838 -514
rect 3342 -1126 3582 -1014
rect 5534 24 5588 514
rect 4094 -566 4920 -514
rect 4094 -1346 4462 -1294
rect 4552 -1346 4920 -1294
rect 5158 -566 5526 -514
rect 5158 -1346 5526 -1294
rect 5536 -2372 5588 -1882
rect 6644 592 6702 692
rect 5748 22 5802 512
rect 6198 -464 6250 24
rect 6644 22 6698 512
rect 7708 592 7766 692
rect 6812 22 6866 512
rect 7262 -464 7314 24
rect 9426 1030 9666 1146
rect 5810 -566 6178 -514
rect 6268 -566 6636 -514
rect 5810 -706 6178 -594
rect 5812 -1126 6180 -1014
rect 5812 -1346 6180 -1294
rect 6270 -1346 6638 -1294
rect 6874 -566 7242 -514
rect 7332 -566 7700 -514
rect 6874 -706 7242 -594
rect 7332 -706 7700 -594
rect 7334 -1126 7702 -1014
rect 6876 -1266 7244 -1154
rect 6876 -1346 7244 -1294
rect 7334 -1346 7702 -1294
rect 5750 -2372 5802 -1882
rect 6200 -1888 6252 -1400
rect 6646 -2372 6700 -1882
rect 5566 -2632 5624 -2532
rect 6814 -2372 6868 -1882
rect 7264 -1882 7316 -1394
rect 6646 -2632 6704 -2532
rect 4478 -2772 4536 -2672
rect 5132 -2912 5190 -2812
rect 7708 -2632 7766 -2532
rect 7260 -2912 7318 -2812
rect 8324 -2772 8382 -2672
rect 3684 -2998 4510 -2946
rect 4748 -2998 5574 -2946
rect 5812 -2998 6180 -2946
rect 6270 -2998 6638 -2946
rect 3542 -5090 3662 -4634
rect 4532 -5090 4726 -4634
rect 6200 -3414 6252 -3038
rect 5596 -5090 5790 -4634
rect 7264 -3414 7316 -3038
rect 8328 -3414 8380 -3038
rect 6876 -3506 7244 -3454
rect 7334 -3506 7702 -3454
rect 6660 -5090 6836 -4634
rect 7940 -3506 8308 -3454
rect 7746 -5090 7896 -4634
<< metal2 >>
rect 3336 3226 9672 3238
rect 3336 2776 3946 3226
rect 4050 2776 4988 3226
rect 5092 2776 5636 3226
rect 5740 2776 6704 3226
rect 6808 2776 7798 3226
rect 7902 2776 9672 3226
rect 3336 2770 9672 2776
rect 8002 1146 9672 1152
rect 8002 1142 9426 1146
rect 8002 1034 8008 1142
rect 8098 1034 9426 1142
rect 8002 1030 9426 1034
rect 9666 1030 9672 1146
rect 8002 1024 9672 1030
rect 5566 692 7766 698
rect 5624 592 6644 692
rect 6702 592 7708 692
rect 5566 586 7766 592
rect 5534 518 5588 520
rect 5534 514 5802 518
rect 5588 512 5802 514
rect 5588 24 5748 512
rect 5534 22 5748 24
rect 6644 512 6866 518
rect 5534 18 5802 22
rect 5748 16 5802 18
rect 6196 24 6252 34
rect 6698 22 6812 512
rect 6644 16 6866 22
rect 7260 24 7316 34
rect 6196 -474 6252 -464
rect 7260 -474 7316 -464
rect 3740 -566 3746 -514
rect 3838 -566 4094 -514
rect 4920 -566 5158 -514
rect 5526 -566 5532 -514
rect 5804 -566 5810 -514
rect 6178 -566 6268 -514
rect 6636 -566 6642 -514
rect 6868 -566 6874 -514
rect 7242 -566 7332 -514
rect 7700 -566 7706 -514
rect 3336 -706 3342 -594
rect 3582 -706 5810 -594
rect 6178 -706 6874 -594
rect 7242 -706 7248 -594
rect 7326 -706 7332 -594
rect 7700 -706 7706 -594
rect 6340 -766 6416 -760
rect 6340 -822 6350 -766
rect 6406 -822 7258 -766
rect 7314 -822 7324 -766
rect 6190 -954 6200 -898
rect 6256 -954 7258 -898
rect 7314 -954 7324 -898
rect 3336 -1126 3342 -1014
rect 3582 -1126 5812 -1014
rect 6180 -1126 7334 -1014
rect 7702 -1126 7708 -1014
rect 6192 -1264 6202 -1208
rect 6258 -1264 6342 -1208
rect 6398 -1264 6408 -1208
rect 6870 -1266 6876 -1154
rect 7244 -1266 7250 -1154
rect 4088 -1346 4094 -1294
rect 4462 -1346 4552 -1294
rect 4920 -1346 5158 -1294
rect 5526 -1346 5532 -1294
rect 5806 -1346 5812 -1294
rect 6180 -1346 6270 -1294
rect 6638 -1346 6644 -1294
rect 6870 -1346 6876 -1294
rect 7244 -1346 7334 -1294
rect 7702 -1346 7708 -1294
rect 6198 -1400 6254 -1390
rect 5536 -1882 5802 -1876
rect 5588 -2372 5750 -1882
rect 7262 -1394 7318 -1384
rect 6198 -1898 6254 -1888
rect 6646 -1882 6868 -1876
rect 5536 -2378 5802 -2372
rect 6700 -2372 6814 -1882
rect 7262 -1892 7318 -1882
rect 6646 -2378 6868 -2372
rect 5566 -2532 7766 -2526
rect 5624 -2632 6646 -2532
rect 6704 -2632 7708 -2532
rect 5566 -2638 7766 -2632
rect 4478 -2668 8382 -2666
rect 4478 -2672 8004 -2668
rect 4536 -2772 8004 -2672
rect 4478 -2776 8004 -2772
rect 8094 -2672 8382 -2668
rect 8094 -2772 8324 -2672
rect 8094 -2776 8382 -2772
rect 4478 -2778 8382 -2776
rect 5132 -2812 7318 -2806
rect 5190 -2912 7260 -2812
rect 5132 -2918 7318 -2912
rect 3678 -2998 3684 -2946
rect 4510 -2998 4516 -2946
rect 4742 -2998 4748 -2946
rect 5574 -2998 5812 -2946
rect 6180 -2998 6270 -2946
rect 6638 -2998 6644 -2946
rect 6198 -3038 6254 -3028
rect 6198 -3454 6254 -3414
rect 7264 -3038 8380 -3032
rect 7316 -3414 8328 -3038
rect 7264 -3420 8380 -3414
rect 8684 -3440 8796 -3414
rect 8684 -3454 8690 -3440
rect 6198 -3506 6876 -3454
rect 7244 -3506 7334 -3454
rect 7702 -3506 7940 -3454
rect 8308 -3504 8690 -3454
rect 8786 -3504 8796 -3440
rect 8308 -3506 8796 -3504
rect 3336 -4634 9672 -4628
rect 3336 -5090 3542 -4634
rect 3662 -5090 4532 -4634
rect 4726 -5090 5596 -4634
rect 5790 -5090 6660 -4634
rect 6836 -5090 7746 -4634
rect 7896 -5090 9672 -4634
rect 3336 -5096 9672 -5090
<< via2 >>
rect 8008 1034 8098 1142
rect 6196 -464 6198 24
rect 6198 -464 6250 24
rect 6250 -464 6252 24
rect 7260 -464 7262 24
rect 7262 -464 7314 24
rect 7314 -464 7316 24
rect 6350 -822 6406 -766
rect 7258 -822 7314 -766
rect 6200 -954 6256 -898
rect 7258 -954 7314 -898
rect 6202 -1264 6258 -1208
rect 6342 -1264 6398 -1208
rect 6198 -1888 6200 -1400
rect 6200 -1888 6252 -1400
rect 6252 -1888 6254 -1400
rect 7262 -1882 7264 -1394
rect 7264 -1882 7316 -1394
rect 7316 -1882 7318 -1394
rect 8004 -2776 8094 -2668
rect 6198 -3414 6200 -3038
rect 6200 -3414 6252 -3038
rect 6252 -3414 6254 -3038
rect 8690 -3504 8786 -3440
<< metal3 >>
rect 8002 1142 8104 1148
rect 8002 1034 8008 1142
rect 8098 1034 8104 1142
rect 8002 1028 8104 1034
rect 6190 24 6258 30
rect 6190 -464 6196 24
rect 6252 -464 6258 24
rect 6190 -892 6258 -464
rect 7254 24 7322 30
rect 7254 -464 7260 24
rect 7316 -464 7322 24
rect 7254 -760 7322 -464
rect 6340 -766 6416 -760
rect 6340 -822 6350 -766
rect 6406 -822 6416 -766
rect 6340 -828 6416 -822
rect 7248 -766 7324 -760
rect 7248 -822 7258 -766
rect 7314 -822 7324 -766
rect 7248 -828 7324 -822
rect 6190 -898 6266 -892
rect 6190 -954 6200 -898
rect 6256 -954 6266 -898
rect 6190 -960 6266 -954
rect 6340 -1202 6408 -828
rect 7248 -898 7324 -892
rect 7248 -954 7258 -898
rect 7314 -954 7324 -898
rect 7248 -960 7324 -954
rect 6192 -1208 6268 -1202
rect 6192 -1264 6202 -1208
rect 6258 -1264 6268 -1208
rect 6192 -1396 6268 -1264
rect 6332 -1208 6408 -1202
rect 6332 -1264 6342 -1208
rect 6398 -1264 6408 -1208
rect 6332 -1270 6408 -1264
rect 7256 -1394 7324 -960
rect 6192 -1400 6260 -1396
rect 6192 -1888 6198 -1400
rect 6254 -1888 6260 -1400
rect 6192 -3038 6260 -1888
rect 7256 -1882 7262 -1394
rect 7318 -1882 7324 -1394
rect 7256 -1894 7324 -1882
rect 7998 -2668 8100 -2662
rect 7998 -2776 8004 -2668
rect 8094 -2776 8100 -2668
rect 7998 -2782 8100 -2776
rect 6192 -3414 6198 -3038
rect 6254 -3414 6260 -3038
rect 6192 -3420 6260 -3414
rect 8684 -3440 8792 -3414
rect 8684 -3504 8690 -3440
rect 8786 -3504 8792 -3440
rect 8684 -3510 8792 -3504
<< via3 >>
rect 8008 1034 8098 1142
rect 8004 -2776 8094 -2668
rect 8690 -3504 8786 -3440
<< metal4 >>
rect 8006 1146 8104 1148
rect 8002 1142 8104 1146
rect 8002 1034 8008 1142
rect 8098 1034 8104 1142
rect 8002 1028 8104 1034
rect 8002 -1376 8098 1028
rect 8002 -2668 8098 -2420
rect 8002 -2776 8004 -2668
rect 8094 -2776 8098 -2668
rect 8002 -2778 8098 -2776
rect 8688 -3440 8788 -2320
rect 8688 -3504 8690 -3440
rect 8786 -3504 8788 -3440
rect 8688 -3506 8788 -3504
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M11
timestamp 1681402674
transform 1 0 5342 0 1 -12
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M12
timestamp 1681402674
transform 1 0 5342 0 1 -1848
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M21
timestamp 1681402674
transform 1 0 5994 0 1 -12
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M22
timestamp 1681402674
transform -1 0 6452 0 1 -12
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M23
timestamp 1681402674
transform -1 0 7518 0 1 -1848
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M24
timestamp 1681402674
transform 1 0 7060 0 1 -1848
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M31
timestamp 1681402674
transform 1 0 7058 0 1 -12
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M32
timestamp 1681402674
transform -1 0 7516 0 1 -12
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M33
timestamp 1681402674
transform -1 0 6454 0 1 -1848
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M34
timestamp 1681402674
transform 1 0 5996 0 1 -1848
box -294 -598 294 564
use sky130_fd_pr__nfet_01v8_lvt_N3YEWU  M41
timestamp 1681226341
transform 1 0 4932 0 1 -3195
box -258 -257 258 257
use sky130_fd_pr__nfet_01v8_lvt_N3YEWU  M42
timestamp 1681226341
transform 1 0 5390 0 1 -3195
box -258 -257 258 257
use sky130_fd_pr__nfet_01v8_lvt_N3YEWU  M51
timestamp 1681226341
transform 1 0 5996 0 1 -3195
box -258 -257 258 257
use sky130_fd_pr__nfet_01v8_lvt_N3YEWU  M52
timestamp 1681226341
transform 1 0 6454 0 1 -3195
box -258 -257 258 257
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M61
timestamp 1681402674
transform -1 0 4736 0 1 -1848
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M62
timestamp 1681402674
transform 1 0 4278 0 1 -1848
box -294 -598 294 564
use sky130_fd_pr__nfet_01v8_lvt_T4X5QS  M71
timestamp 1681226341
transform 1 0 7060 0 1 -3257
box -258 -257 258 257
use sky130_fd_pr__nfet_01v8_lvt_T4X5QS  M72
timestamp 1681226341
transform 1 0 7518 0 1 -3257
box -258 -257 258 257
use sky130_fd_pr__nfet_01v8_lvt_T4X5QS  M73
timestamp 1681226341
transform 1 0 8124 0 1 -3257
box -258 -257 258 257
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M81
timestamp 1681402674
transform 1 0 4278 0 1 -12
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M82
timestamp 1681402674
transform -1 0 4736 0 1 -12
box -294 -564 294 598
use sky130_fd_pr__nfet_01v8_lvt_N3YEWU  M91
timestamp 1681226341
transform 1 0 3868 0 1 -3195
box -258 -257 258 257
use sky130_fd_pr__nfet_01v8_lvt_N3YEWU  M92
timestamp 1681226341
transform -1 0 4326 0 1 -3195
box -258 -257 258 257
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  XC2
timestamp 1680255405
transform -1 0 8684 0 1 -1900
box -686 -540 686 540
<< labels >>
flabel metal1 3336 -2262 3588 -968 0 FreeMono 1280 90 0 0 vinp
port 2 nsew
flabel metal1 3336 -752 3588 542 0 FreeMono 1280 90 0 0 vinn
port 3 nsew
flabel metal2 3336 2770 9672 3238 0 FreeMono 1280 0 0 0 vdd
port 0 nsew
flabel metal2 3336 -5096 9672 -4628 0 FreeMono 1280 0 0 0 vss
port 1 nsew
flabel metal1 9420 836 9672 2130 0 FreeMono 1280 90 0 0 out
port 4 nsew
<< end >>
