magic
tech sky130A
magscale 1 2
timestamp 1680252321
<< xpolycontact >>
rect -35 350 35 782
rect -35 -782 35 -350
<< xpolyres >>
rect -35 -350 35 350
<< viali >>
rect -19 367 19 764
rect -19 -764 19 -367
<< metal1 >>
rect -25 764 25 776
rect -25 367 -19 764
rect 19 367 25 764
rect -25 355 25 367
rect -25 -367 25 -355
rect -25 -764 -19 -367
rect 19 -764 25 -367
rect -25 -776 25 -764
<< res0p35 >>
rect -37 -352 37 352
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 3.5 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 21.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
