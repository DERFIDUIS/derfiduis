** sch_path:
*+ /home/antony/Documentos/Xschem-Projects/WORK_IN_PROGRESS/My_xschem/For_Layout/BGR_lvt.sch
.subckt BGR_lvt vdd vss out
*.PININFO vdd:B vss:B out:B
M1 net3 net3 net5 vss sky130_fd_pr__nfet_01v8_lvt L=7 W=5 nf=1 m=1
M2 net5 net5 vss vss sky130_fd_pr__nfet_01v8_lvt L=7 W=5 nf=1 m=1
M31 net3 net2 net1 vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 m=1
M41 net1 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 m=1
M51 net4 net3 net2 vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 m=1
M61 net4 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M71 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M81 net4 net4 net6 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M91 net2 net4 net8 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
Q1 vss vss net6 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
Q21 vss vss net7 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
M101 out net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
Q3 vss vss net9 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
XR3 net7 net8 vss sky130_fd_pr__res_xhigh_po_0p69 L=0.94 mult=1 m=1
XR4 net9 out vss sky130_fd_pr__res_xhigh_po_0p69 L=6 mult=1 m=1
M42 net1 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 m=1
M32 net3 net2 net1 vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=5 nf=1 m=1
M52 net4 net3 net2 vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=2 nf=1 m=1
M62 net4 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M63 net4 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M64 net4 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M65 net4 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M66 net4 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M82 net4 net4 net6 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M83 net4 net4 net6 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M84 net4 net4 net6 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M85 net4 net4 net6 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M86 net4 net4 net6 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M72 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M73 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M74 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M75 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M76 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M92 net2 net4 net8 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M93 net2 net4 net8 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M94 net2 net4 net8 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M95 net2 net4 net8 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M96 net2 net4 net8 vss sky130_fd_pr__nfet_01v8_lvt L=2 W=5 nf=1 m=1
M102 out net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M103 out net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M104 out net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M105 out net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M106 out net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
Q22 vss vss net7 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
Q23 vss vss net7 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
Q24 vss vss net7 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
Q25 vss vss net7 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
Q26 vss vss net7 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
Q27 vss vss net7 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
Q28 vss vss net7 sky130_fd_pr__pnp_05v5_W3p40L3p40 NE=1 m=1
.ends
.end
