magic
tech sky130A
magscale 1 2
timestamp 1680265380
<< error_p >>
rect -31 581 31 587
rect -31 547 -19 581
rect -31 541 31 547
rect -31 -547 31 -541
rect -31 -581 -19 -547
rect -31 -587 31 -581
<< nwell >>
rect -231 -719 231 719
<< pmoslvt >>
rect -35 -500 35 500
<< pdiff >>
rect -93 488 -35 500
rect -93 -488 -81 488
rect -47 -488 -35 488
rect -93 -500 -35 -488
rect 35 488 93 500
rect 35 -488 47 488
rect 81 -488 93 488
rect 35 -500 93 -488
<< pdiffc >>
rect -81 -488 -47 488
rect 47 -488 81 488
<< nsubdiff >>
rect -195 649 -99 683
rect 99 649 195 683
rect -195 587 -161 649
rect 161 587 195 649
rect -195 -649 -161 -587
rect 161 -649 195 -587
rect -195 -683 -99 -649
rect 99 -683 195 -649
<< nsubdiffcont >>
rect -99 649 99 683
rect -195 -587 -161 587
rect 161 -587 195 587
rect -99 -683 99 -649
<< poly >>
rect -35 581 35 597
rect -35 547 -19 581
rect 19 547 35 581
rect -35 500 35 547
rect -35 -547 35 -500
rect -35 -581 -19 -547
rect 19 -581 35 -547
rect -35 -597 35 -581
<< polycont >>
rect -19 547 19 581
rect -19 -581 19 -547
<< locali >>
rect -195 649 -99 683
rect 99 649 195 683
rect -195 587 -161 649
rect 161 587 195 649
rect -35 547 -19 581
rect 19 547 35 581
rect -81 488 -47 504
rect -81 -504 -47 -488
rect 47 488 81 504
rect 47 -504 81 -488
rect -35 -581 -19 -547
rect 19 -581 35 -547
rect -195 -649 -161 -587
rect 161 -649 195 -587
rect -195 -683 -99 -649
rect 99 -683 195 -649
<< viali >>
rect -19 547 19 581
rect -81 -488 -47 488
rect 47 -488 81 488
rect -19 -581 19 -547
<< metal1 >>
rect -31 581 31 587
rect -31 547 -19 581
rect 19 547 31 581
rect -31 541 31 547
rect -87 488 -41 500
rect -87 -488 -81 488
rect -47 -488 -41 488
rect -87 -500 -41 -488
rect 41 488 87 500
rect 41 -488 47 488
rect 81 -488 87 488
rect 41 -500 87 -488
rect -31 -547 31 -541
rect -31 -581 -19 -547
rect 19 -581 31 -547
rect -31 -587 31 -581
<< properties >>
string FIXED_BBOX -178 -666 178 666
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
