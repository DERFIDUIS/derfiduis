magic
tech sky130A
magscale 1 2
timestamp 1681878372
<< nwell >>
rect 2002 -3900 2068 -2738
rect 2402 -3900 2516 -2738
rect 3472 -3900 3586 -2738
rect 4536 -3900 4650 -2738
rect 5600 -3900 5714 -2738
rect 6664 -3900 6778 -2738
rect 7906 -3460 7972 -3336
rect 7898 -3494 7972 -3460
rect 7906 -3532 7972 -3494
rect 7898 -3566 7972 -3532
rect 7906 -3600 7972 -3566
rect 7898 -3634 7972 -3600
rect 7906 -3668 7972 -3634
rect 7898 -3702 7972 -3668
rect 7906 -3898 7972 -3702
rect 2002 -5448 2068 -4286
rect 2408 -5448 2522 -4286
rect 3472 -5448 3586 -4286
rect 4536 -5448 4650 -4286
rect 5600 -5448 5714 -4286
rect 6664 -5448 6778 -4286
rect 7806 -4348 7864 -4344
rect 7906 -4448 7972 -4286
rect 7898 -4482 7972 -4448
rect 7906 -4520 7972 -4482
rect 7898 -4554 7972 -4520
rect 7906 -4588 7972 -4554
rect 7898 -4622 7972 -4588
rect 7906 -4656 7972 -4622
rect 7898 -4690 7972 -4656
rect 7906 -4848 7972 -4690
<< pwell >>
rect 1146 -8312 1384 -7260
rect 8938 -7950 9174 -5886
<< nbase >>
rect 3796 -8868 3858 -8578
rect 4612 -8868 4674 -8578
rect 5428 -8868 5490 -8578
rect 6244 -8868 6306 -8578
rect 7060 -8868 7122 -8578
rect 3796 -9684 3858 -9394
rect 4612 -9684 4674 -9394
rect 5428 -9684 5490 -9394
rect 6244 -9684 6306 -9394
rect 7060 -9684 7122 -9394
<< ndiff >>
rect 9556 -4248 9558 -3248
rect 9556 -5404 9558 -4404
rect 1702 -7146 1704 -6146
rect 2678 -7146 2680 -6146
rect 2766 -7146 2768 -6146
rect 3742 -7146 3744 -6146
rect 3830 -7146 3832 -6146
rect 4806 -7146 4808 -6146
rect 5966 -7146 5968 -6146
rect 6054 -7146 6056 -6146
rect 7030 -7146 7032 -6146
rect 7118 -7146 7120 -6146
rect 8094 -7146 8096 -6146
rect 8182 -7146 8184 -6146
<< pdiff >>
rect 1966 -3800 1968 -2800
rect 2420 -3800 2422 -2800
rect 2508 -3800 2510 -2800
rect 3484 -3800 3486 -2800
rect 3572 -3800 3574 -2800
rect 4548 -3800 4550 -2800
rect 4636 -3800 4638 -2800
rect 5612 -3800 5614 -2800
rect 5700 -3800 5702 -2800
rect 6676 -3800 6678 -2800
rect 6764 -3800 6766 -2800
rect 7870 -3798 7872 -3398
rect 1966 -5386 1968 -4386
rect 2420 -5386 2422 -4386
rect 2508 -5386 2510 -4386
rect 3484 -5386 3486 -4386
rect 3572 -5386 3574 -4386
rect 4548 -5386 4550 -4386
rect 4636 -5386 4638 -4386
rect 5612 -5386 5614 -4386
rect 5700 -5386 5702 -4386
rect 6676 -5386 6678 -4386
rect 6764 -5386 6766 -4386
rect 7870 -4786 7872 -4386
<< psubdiff >>
rect 9558 -3302 9622 -3248
rect 9558 -3336 9584 -3302
rect 9618 -3336 9622 -3302
rect 9558 -3370 9622 -3336
rect 9558 -3404 9584 -3370
rect 9618 -3404 9622 -3370
rect 9558 -3438 9622 -3404
rect 9558 -3472 9584 -3438
rect 9618 -3472 9622 -3438
rect 9558 -3506 9622 -3472
rect 9558 -3540 9584 -3506
rect 9618 -3540 9622 -3506
rect 9558 -3574 9622 -3540
rect 9558 -3608 9584 -3574
rect 9618 -3608 9622 -3574
rect 9558 -3642 9622 -3608
rect 9558 -3676 9584 -3642
rect 9618 -3676 9622 -3642
rect 9558 -3710 9622 -3676
rect 9558 -3744 9584 -3710
rect 9618 -3744 9622 -3710
rect 9558 -3778 9622 -3744
rect 9558 -3812 9584 -3778
rect 9618 -3812 9622 -3778
rect 9558 -3846 9622 -3812
rect 9558 -3880 9584 -3846
rect 9618 -3880 9622 -3846
rect 9558 -3914 9622 -3880
rect 9558 -3948 9584 -3914
rect 9618 -3948 9622 -3914
rect 9558 -3982 9622 -3948
rect 9558 -4016 9584 -3982
rect 9618 -4016 9622 -3982
rect 9558 -4050 9622 -4016
rect 9558 -4084 9584 -4050
rect 9618 -4084 9622 -4050
rect 9558 -4118 9622 -4084
rect 9558 -4152 9584 -4118
rect 9618 -4152 9622 -4118
rect 9558 -4186 9622 -4152
rect 9558 -4220 9584 -4186
rect 9618 -4220 9622 -4186
rect 9558 -4248 9622 -4220
rect 9558 -4458 9622 -4404
rect 9558 -4492 9584 -4458
rect 9618 -4492 9622 -4458
rect 9558 -4526 9622 -4492
rect 9558 -4560 9584 -4526
rect 9618 -4560 9622 -4526
rect 9558 -4594 9622 -4560
rect 9558 -4628 9584 -4594
rect 9618 -4628 9622 -4594
rect 9558 -4662 9622 -4628
rect 9558 -4696 9584 -4662
rect 9618 -4696 9622 -4662
rect 9558 -4730 9622 -4696
rect 9558 -4764 9584 -4730
rect 9618 -4764 9622 -4730
rect 9558 -4798 9622 -4764
rect 9558 -4832 9584 -4798
rect 9618 -4832 9622 -4798
rect 9558 -4866 9622 -4832
rect 9558 -4900 9584 -4866
rect 9618 -4900 9622 -4866
rect 9558 -4934 9622 -4900
rect 9558 -4968 9584 -4934
rect 9618 -4968 9622 -4934
rect 9558 -5002 9622 -4968
rect 9558 -5036 9584 -5002
rect 9618 -5036 9622 -5002
rect 9558 -5070 9622 -5036
rect 9558 -5104 9584 -5070
rect 9618 -5104 9622 -5070
rect 9558 -5138 9622 -5104
rect 9558 -5172 9584 -5138
rect 9618 -5172 9622 -5138
rect 9558 -5206 9622 -5172
rect 9558 -5240 9584 -5206
rect 9618 -5240 9622 -5206
rect 9558 -5274 9622 -5240
rect 9558 -5308 9584 -5274
rect 9618 -5308 9622 -5274
rect 9558 -5342 9622 -5308
rect 9558 -5376 9584 -5342
rect 9618 -5376 9622 -5342
rect 9558 -5404 9622 -5376
rect 8938 -5978 9066 -5886
rect 1638 -6200 1702 -6146
rect 1638 -6234 1642 -6200
rect 1676 -6234 1702 -6200
rect 1638 -6268 1702 -6234
rect 1638 -6302 1642 -6268
rect 1676 -6302 1702 -6268
rect 1638 -6336 1702 -6302
rect 1638 -6370 1642 -6336
rect 1676 -6370 1702 -6336
rect 1638 -6404 1702 -6370
rect 1638 -6438 1642 -6404
rect 1676 -6438 1702 -6404
rect 1638 -6472 1702 -6438
rect 1638 -6506 1642 -6472
rect 1676 -6506 1702 -6472
rect 1638 -6540 1702 -6506
rect 1638 -6574 1642 -6540
rect 1676 -6574 1702 -6540
rect 1638 -6608 1702 -6574
rect 1638 -6642 1642 -6608
rect 1676 -6642 1702 -6608
rect 1638 -6676 1702 -6642
rect 1638 -6710 1642 -6676
rect 1676 -6710 1702 -6676
rect 1638 -6744 1702 -6710
rect 1638 -6778 1642 -6744
rect 1676 -6778 1702 -6744
rect 1638 -6812 1702 -6778
rect 1638 -6846 1642 -6812
rect 1676 -6846 1702 -6812
rect 1638 -6880 1702 -6846
rect 1638 -6914 1642 -6880
rect 1676 -6914 1702 -6880
rect 1638 -6948 1702 -6914
rect 1638 -6982 1642 -6948
rect 1676 -6982 1702 -6948
rect 1638 -7016 1702 -6982
rect 1638 -7050 1642 -7016
rect 1676 -7050 1702 -7016
rect 1638 -7084 1702 -7050
rect 1638 -7118 1642 -7084
rect 1676 -7118 1702 -7084
rect 1638 -7146 1702 -7118
rect 2680 -6200 2766 -6146
rect 2680 -6234 2706 -6200
rect 2740 -6234 2766 -6200
rect 2680 -6268 2766 -6234
rect 2680 -6302 2706 -6268
rect 2740 -6302 2766 -6268
rect 2680 -6336 2766 -6302
rect 2680 -6370 2706 -6336
rect 2740 -6370 2766 -6336
rect 2680 -6404 2766 -6370
rect 2680 -6438 2706 -6404
rect 2740 -6438 2766 -6404
rect 2680 -6472 2766 -6438
rect 2680 -6506 2706 -6472
rect 2740 -6506 2766 -6472
rect 2680 -6540 2766 -6506
rect 2680 -6574 2706 -6540
rect 2740 -6574 2766 -6540
rect 2680 -6608 2766 -6574
rect 2680 -6642 2706 -6608
rect 2740 -6642 2766 -6608
rect 2680 -6676 2766 -6642
rect 2680 -6710 2706 -6676
rect 2740 -6710 2766 -6676
rect 2680 -6744 2766 -6710
rect 2680 -6778 2706 -6744
rect 2740 -6778 2766 -6744
rect 2680 -6812 2766 -6778
rect 2680 -6846 2706 -6812
rect 2740 -6846 2766 -6812
rect 2680 -6880 2766 -6846
rect 2680 -6914 2706 -6880
rect 2740 -6914 2766 -6880
rect 2680 -6948 2766 -6914
rect 2680 -6982 2706 -6948
rect 2740 -6982 2766 -6948
rect 2680 -7016 2766 -6982
rect 2680 -7050 2706 -7016
rect 2740 -7050 2766 -7016
rect 2680 -7084 2766 -7050
rect 2680 -7118 2706 -7084
rect 2740 -7118 2766 -7084
rect 2680 -7146 2766 -7118
rect 3744 -6200 3830 -6146
rect 3744 -6234 3770 -6200
rect 3804 -6234 3830 -6200
rect 3744 -6268 3830 -6234
rect 3744 -6302 3770 -6268
rect 3804 -6302 3830 -6268
rect 3744 -6336 3830 -6302
rect 3744 -6370 3770 -6336
rect 3804 -6370 3830 -6336
rect 3744 -6404 3830 -6370
rect 3744 -6438 3770 -6404
rect 3804 -6438 3830 -6404
rect 3744 -6472 3830 -6438
rect 3744 -6506 3770 -6472
rect 3804 -6506 3830 -6472
rect 3744 -6540 3830 -6506
rect 3744 -6574 3770 -6540
rect 3804 -6574 3830 -6540
rect 3744 -6608 3830 -6574
rect 3744 -6642 3770 -6608
rect 3804 -6642 3830 -6608
rect 3744 -6676 3830 -6642
rect 3744 -6710 3770 -6676
rect 3804 -6710 3830 -6676
rect 3744 -6744 3830 -6710
rect 3744 -6778 3770 -6744
rect 3804 -6778 3830 -6744
rect 3744 -6812 3830 -6778
rect 3744 -6846 3770 -6812
rect 3804 -6846 3830 -6812
rect 3744 -6880 3830 -6846
rect 3744 -6914 3770 -6880
rect 3804 -6914 3830 -6880
rect 3744 -6948 3830 -6914
rect 3744 -6982 3770 -6948
rect 3804 -6982 3830 -6948
rect 3744 -7016 3830 -6982
rect 3744 -7050 3770 -7016
rect 3804 -7050 3830 -7016
rect 3744 -7084 3830 -7050
rect 3744 -7118 3770 -7084
rect 3804 -7118 3830 -7084
rect 3744 -7146 3830 -7118
rect 4808 -6200 4872 -6146
rect 4808 -6234 4834 -6200
rect 4868 -6234 4872 -6200
rect 4808 -6268 4872 -6234
rect 4808 -6302 4834 -6268
rect 4868 -6302 4872 -6268
rect 4808 -6336 4872 -6302
rect 4808 -6370 4834 -6336
rect 4868 -6370 4872 -6336
rect 4808 -6404 4872 -6370
rect 4808 -6438 4834 -6404
rect 4868 -6438 4872 -6404
rect 4808 -6472 4872 -6438
rect 4808 -6506 4834 -6472
rect 4868 -6506 4872 -6472
rect 4808 -6540 4872 -6506
rect 4808 -6574 4834 -6540
rect 4868 -6574 4872 -6540
rect 4808 -6608 4872 -6574
rect 4808 -6642 4834 -6608
rect 4868 -6642 4872 -6608
rect 4808 -6676 4872 -6642
rect 4808 -6710 4834 -6676
rect 4868 -6710 4872 -6676
rect 4808 -6744 4872 -6710
rect 4808 -6778 4834 -6744
rect 4868 -6778 4872 -6744
rect 4808 -6812 4872 -6778
rect 4808 -6846 4834 -6812
rect 4868 -6846 4872 -6812
rect 4808 -6880 4872 -6846
rect 4808 -6914 4834 -6880
rect 4868 -6914 4872 -6880
rect 4808 -6948 4872 -6914
rect 4808 -6982 4834 -6948
rect 4868 -6982 4872 -6948
rect 4808 -7016 4872 -6982
rect 4808 -7050 4834 -7016
rect 4868 -7050 4872 -7016
rect 4808 -7084 4872 -7050
rect 4808 -7118 4834 -7084
rect 4868 -7118 4872 -7084
rect 4808 -7146 4872 -7118
rect 5968 -6200 6054 -6146
rect 5968 -6234 5994 -6200
rect 6028 -6234 6054 -6200
rect 5968 -6268 6054 -6234
rect 5968 -6302 5994 -6268
rect 6028 -6302 6054 -6268
rect 5968 -6336 6054 -6302
rect 5968 -6370 5994 -6336
rect 6028 -6370 6054 -6336
rect 5968 -6404 6054 -6370
rect 5968 -6438 5994 -6404
rect 6028 -6438 6054 -6404
rect 5968 -6472 6054 -6438
rect 5968 -6506 5994 -6472
rect 6028 -6506 6054 -6472
rect 5968 -6540 6054 -6506
rect 5968 -6574 5994 -6540
rect 6028 -6574 6054 -6540
rect 5968 -6608 6054 -6574
rect 5968 -6642 5994 -6608
rect 6028 -6642 6054 -6608
rect 5968 -6676 6054 -6642
rect 5968 -6710 5994 -6676
rect 6028 -6710 6054 -6676
rect 5968 -6744 6054 -6710
rect 5968 -6778 5994 -6744
rect 6028 -6778 6054 -6744
rect 5968 -6812 6054 -6778
rect 5968 -6846 5994 -6812
rect 6028 -6846 6054 -6812
rect 5968 -6880 6054 -6846
rect 5968 -6914 5994 -6880
rect 6028 -6914 6054 -6880
rect 5968 -6948 6054 -6914
rect 5968 -6982 5994 -6948
rect 6028 -6982 6054 -6948
rect 5968 -7016 6054 -6982
rect 5968 -7050 5994 -7016
rect 6028 -7050 6054 -7016
rect 5968 -7084 6054 -7050
rect 5968 -7118 5994 -7084
rect 6028 -7118 6054 -7084
rect 5968 -7146 6054 -7118
rect 7032 -6200 7118 -6146
rect 7032 -6234 7058 -6200
rect 7092 -6234 7118 -6200
rect 7032 -6268 7118 -6234
rect 7032 -6302 7058 -6268
rect 7092 -6302 7118 -6268
rect 7032 -6336 7118 -6302
rect 7032 -6370 7058 -6336
rect 7092 -6370 7118 -6336
rect 7032 -6404 7118 -6370
rect 7032 -6438 7058 -6404
rect 7092 -6438 7118 -6404
rect 7032 -6472 7118 -6438
rect 7032 -6506 7058 -6472
rect 7092 -6506 7118 -6472
rect 7032 -6540 7118 -6506
rect 7032 -6574 7058 -6540
rect 7092 -6574 7118 -6540
rect 7032 -6608 7118 -6574
rect 7032 -6642 7058 -6608
rect 7092 -6642 7118 -6608
rect 7032 -6676 7118 -6642
rect 7032 -6710 7058 -6676
rect 7092 -6710 7118 -6676
rect 7032 -6744 7118 -6710
rect 7032 -6778 7058 -6744
rect 7092 -6778 7118 -6744
rect 7032 -6812 7118 -6778
rect 7032 -6846 7058 -6812
rect 7092 -6846 7118 -6812
rect 7032 -6880 7118 -6846
rect 7032 -6914 7058 -6880
rect 7092 -6914 7118 -6880
rect 7032 -6948 7118 -6914
rect 7032 -6982 7058 -6948
rect 7092 -6982 7118 -6948
rect 7032 -7016 7118 -6982
rect 7032 -7050 7058 -7016
rect 7092 -7050 7118 -7016
rect 7032 -7084 7118 -7050
rect 7032 -7118 7058 -7084
rect 7092 -7118 7118 -7084
rect 7032 -7146 7118 -7118
rect 8096 -6200 8182 -6146
rect 8096 -6234 8122 -6200
rect 8156 -6234 8182 -6200
rect 8096 -6268 8182 -6234
rect 8096 -6302 8122 -6268
rect 8156 -6302 8182 -6268
rect 8096 -6336 8182 -6302
rect 8096 -6370 8122 -6336
rect 8156 -6370 8182 -6336
rect 8096 -6404 8182 -6370
rect 8096 -6438 8122 -6404
rect 8156 -6438 8182 -6404
rect 8096 -6472 8182 -6438
rect 8096 -6506 8122 -6472
rect 8156 -6506 8182 -6472
rect 8096 -6540 8182 -6506
rect 8096 -6574 8122 -6540
rect 8156 -6574 8182 -6540
rect 8096 -6608 8182 -6574
rect 8096 -6642 8122 -6608
rect 8156 -6642 8182 -6608
rect 8096 -6676 8182 -6642
rect 8096 -6710 8122 -6676
rect 8156 -6710 8182 -6676
rect 8096 -6744 8182 -6710
rect 8096 -6778 8122 -6744
rect 8156 -6778 8182 -6744
rect 8096 -6812 8182 -6778
rect 8096 -6846 8122 -6812
rect 8156 -6846 8182 -6812
rect 8096 -6880 8182 -6846
rect 8096 -6914 8122 -6880
rect 8156 -6914 8182 -6880
rect 8096 -6948 8182 -6914
rect 8096 -6982 8122 -6948
rect 8156 -6982 8182 -6948
rect 8096 -7016 8182 -6982
rect 8096 -7050 8122 -7016
rect 8156 -7050 8182 -7016
rect 8096 -7084 8182 -7050
rect 8096 -7118 8122 -7084
rect 8156 -7118 8182 -7084
rect 8096 -7146 8182 -7118
rect 8938 -6150 8962 -5978
rect 9042 -6150 9066 -5978
rect 8938 -6322 9066 -6150
rect 8938 -6494 8962 -6322
rect 9042 -6494 9066 -6322
rect 8938 -6666 9066 -6494
rect 8938 -6838 8962 -6666
rect 9042 -6838 9066 -6666
rect 8938 -7010 9066 -6838
rect 8938 -7182 8962 -7010
rect 9042 -7182 9066 -7010
rect 1146 -7418 1274 -7260
rect 1146 -7590 1170 -7418
rect 1250 -7590 1274 -7418
rect 1146 -7762 1274 -7590
rect 1146 -7934 1170 -7762
rect 1250 -7934 1274 -7762
rect 1146 -8106 1274 -7934
rect 8938 -7354 9066 -7182
rect 8938 -7526 8962 -7354
rect 9042 -7526 9066 -7354
rect 8938 -7698 9066 -7526
rect 8938 -7870 8962 -7698
rect 9042 -7870 9066 -7698
rect 8938 -7950 9066 -7870
rect 1146 -8278 1170 -8106
rect 1250 -8278 1274 -8106
rect 1146 -8312 1274 -8278
<< nsubdiff >>
rect 1968 -2854 2032 -2800
rect 1968 -2888 1994 -2854
rect 2028 -2888 2032 -2854
rect 1968 -2922 2032 -2888
rect 1968 -2956 1994 -2922
rect 2028 -2956 2032 -2922
rect 1968 -2990 2032 -2956
rect 1968 -3024 1994 -2990
rect 2028 -3024 2032 -2990
rect 1968 -3058 2032 -3024
rect 1968 -3092 1994 -3058
rect 2028 -3092 2032 -3058
rect 1968 -3126 2032 -3092
rect 1968 -3160 1994 -3126
rect 2028 -3160 2032 -3126
rect 1968 -3194 2032 -3160
rect 1968 -3228 1994 -3194
rect 2028 -3228 2032 -3194
rect 1968 -3262 2032 -3228
rect 1968 -3296 1994 -3262
rect 2028 -3296 2032 -3262
rect 1968 -3330 2032 -3296
rect 1968 -3364 1994 -3330
rect 2028 -3364 2032 -3330
rect 1968 -3398 2032 -3364
rect 1968 -3432 1994 -3398
rect 2028 -3432 2032 -3398
rect 1968 -3466 2032 -3432
rect 1968 -3500 1994 -3466
rect 2028 -3500 2032 -3466
rect 1968 -3534 2032 -3500
rect 1968 -3568 1994 -3534
rect 2028 -3568 2032 -3534
rect 1968 -3602 2032 -3568
rect 1968 -3636 1994 -3602
rect 2028 -3636 2032 -3602
rect 1968 -3670 2032 -3636
rect 1968 -3704 1994 -3670
rect 2028 -3704 2032 -3670
rect 1968 -3738 2032 -3704
rect 1968 -3772 1994 -3738
rect 2028 -3772 2032 -3738
rect 1968 -3800 2032 -3772
rect 2422 -2854 2508 -2800
rect 2422 -2888 2448 -2854
rect 2482 -2888 2508 -2854
rect 2422 -2922 2508 -2888
rect 2422 -2956 2448 -2922
rect 2482 -2956 2508 -2922
rect 2422 -2990 2508 -2956
rect 2422 -3024 2448 -2990
rect 2482 -3024 2508 -2990
rect 2422 -3058 2508 -3024
rect 2422 -3092 2448 -3058
rect 2482 -3092 2508 -3058
rect 2422 -3126 2508 -3092
rect 2422 -3160 2448 -3126
rect 2482 -3160 2508 -3126
rect 2422 -3194 2508 -3160
rect 2422 -3228 2448 -3194
rect 2482 -3228 2508 -3194
rect 2422 -3262 2508 -3228
rect 2422 -3296 2448 -3262
rect 2482 -3296 2508 -3262
rect 2422 -3330 2508 -3296
rect 2422 -3364 2448 -3330
rect 2482 -3364 2508 -3330
rect 2422 -3398 2508 -3364
rect 2422 -3432 2448 -3398
rect 2482 -3432 2508 -3398
rect 2422 -3466 2508 -3432
rect 2422 -3500 2448 -3466
rect 2482 -3500 2508 -3466
rect 2422 -3534 2508 -3500
rect 2422 -3568 2448 -3534
rect 2482 -3568 2508 -3534
rect 2422 -3602 2508 -3568
rect 2422 -3636 2448 -3602
rect 2482 -3636 2508 -3602
rect 2422 -3670 2508 -3636
rect 2422 -3704 2448 -3670
rect 2482 -3704 2508 -3670
rect 2422 -3738 2508 -3704
rect 2422 -3772 2448 -3738
rect 2482 -3772 2508 -3738
rect 2422 -3800 2508 -3772
rect 3486 -2854 3572 -2800
rect 3486 -2888 3512 -2854
rect 3546 -2888 3572 -2854
rect 3486 -2922 3572 -2888
rect 3486 -2956 3512 -2922
rect 3546 -2956 3572 -2922
rect 3486 -2990 3572 -2956
rect 3486 -3024 3512 -2990
rect 3546 -3024 3572 -2990
rect 3486 -3058 3572 -3024
rect 3486 -3092 3512 -3058
rect 3546 -3092 3572 -3058
rect 3486 -3126 3572 -3092
rect 3486 -3160 3512 -3126
rect 3546 -3160 3572 -3126
rect 3486 -3194 3572 -3160
rect 3486 -3228 3512 -3194
rect 3546 -3228 3572 -3194
rect 3486 -3262 3572 -3228
rect 3486 -3296 3512 -3262
rect 3546 -3296 3572 -3262
rect 3486 -3330 3572 -3296
rect 3486 -3364 3512 -3330
rect 3546 -3364 3572 -3330
rect 3486 -3398 3572 -3364
rect 3486 -3432 3512 -3398
rect 3546 -3432 3572 -3398
rect 3486 -3466 3572 -3432
rect 3486 -3500 3512 -3466
rect 3546 -3500 3572 -3466
rect 3486 -3534 3572 -3500
rect 3486 -3568 3512 -3534
rect 3546 -3568 3572 -3534
rect 3486 -3602 3572 -3568
rect 3486 -3636 3512 -3602
rect 3546 -3636 3572 -3602
rect 3486 -3670 3572 -3636
rect 3486 -3704 3512 -3670
rect 3546 -3704 3572 -3670
rect 3486 -3738 3572 -3704
rect 3486 -3772 3512 -3738
rect 3546 -3772 3572 -3738
rect 3486 -3800 3572 -3772
rect 4550 -2854 4636 -2800
rect 4550 -2888 4576 -2854
rect 4610 -2888 4636 -2854
rect 4550 -2922 4636 -2888
rect 4550 -2956 4576 -2922
rect 4610 -2956 4636 -2922
rect 4550 -2990 4636 -2956
rect 4550 -3024 4576 -2990
rect 4610 -3024 4636 -2990
rect 4550 -3058 4636 -3024
rect 4550 -3092 4576 -3058
rect 4610 -3092 4636 -3058
rect 4550 -3126 4636 -3092
rect 4550 -3160 4576 -3126
rect 4610 -3160 4636 -3126
rect 4550 -3194 4636 -3160
rect 4550 -3228 4576 -3194
rect 4610 -3228 4636 -3194
rect 4550 -3262 4636 -3228
rect 4550 -3296 4576 -3262
rect 4610 -3296 4636 -3262
rect 4550 -3330 4636 -3296
rect 4550 -3364 4576 -3330
rect 4610 -3364 4636 -3330
rect 4550 -3398 4636 -3364
rect 4550 -3432 4576 -3398
rect 4610 -3432 4636 -3398
rect 4550 -3466 4636 -3432
rect 4550 -3500 4576 -3466
rect 4610 -3500 4636 -3466
rect 4550 -3534 4636 -3500
rect 4550 -3568 4576 -3534
rect 4610 -3568 4636 -3534
rect 4550 -3602 4636 -3568
rect 4550 -3636 4576 -3602
rect 4610 -3636 4636 -3602
rect 4550 -3670 4636 -3636
rect 4550 -3704 4576 -3670
rect 4610 -3704 4636 -3670
rect 4550 -3738 4636 -3704
rect 4550 -3772 4576 -3738
rect 4610 -3772 4636 -3738
rect 4550 -3800 4636 -3772
rect 5614 -2854 5700 -2800
rect 5614 -2888 5640 -2854
rect 5674 -2888 5700 -2854
rect 5614 -2922 5700 -2888
rect 5614 -2956 5640 -2922
rect 5674 -2956 5700 -2922
rect 5614 -2990 5700 -2956
rect 5614 -3024 5640 -2990
rect 5674 -3024 5700 -2990
rect 5614 -3058 5700 -3024
rect 5614 -3092 5640 -3058
rect 5674 -3092 5700 -3058
rect 5614 -3126 5700 -3092
rect 5614 -3160 5640 -3126
rect 5674 -3160 5700 -3126
rect 5614 -3194 5700 -3160
rect 5614 -3228 5640 -3194
rect 5674 -3228 5700 -3194
rect 5614 -3262 5700 -3228
rect 5614 -3296 5640 -3262
rect 5674 -3296 5700 -3262
rect 5614 -3330 5700 -3296
rect 5614 -3364 5640 -3330
rect 5674 -3364 5700 -3330
rect 5614 -3398 5700 -3364
rect 5614 -3432 5640 -3398
rect 5674 -3432 5700 -3398
rect 5614 -3466 5700 -3432
rect 5614 -3500 5640 -3466
rect 5674 -3500 5700 -3466
rect 5614 -3534 5700 -3500
rect 5614 -3568 5640 -3534
rect 5674 -3568 5700 -3534
rect 5614 -3602 5700 -3568
rect 5614 -3636 5640 -3602
rect 5674 -3636 5700 -3602
rect 5614 -3670 5700 -3636
rect 5614 -3704 5640 -3670
rect 5674 -3704 5700 -3670
rect 5614 -3738 5700 -3704
rect 5614 -3772 5640 -3738
rect 5674 -3772 5700 -3738
rect 5614 -3800 5700 -3772
rect 6678 -2854 6764 -2800
rect 6678 -2888 6704 -2854
rect 6738 -2888 6764 -2854
rect 6678 -2922 6764 -2888
rect 6678 -2956 6704 -2922
rect 6738 -2956 6764 -2922
rect 6678 -2990 6764 -2956
rect 6678 -3024 6704 -2990
rect 6738 -3024 6764 -2990
rect 6678 -3058 6764 -3024
rect 6678 -3092 6704 -3058
rect 6738 -3092 6764 -3058
rect 6678 -3126 6764 -3092
rect 6678 -3160 6704 -3126
rect 6738 -3160 6764 -3126
rect 6678 -3194 6764 -3160
rect 6678 -3228 6704 -3194
rect 6738 -3228 6764 -3194
rect 6678 -3262 6764 -3228
rect 6678 -3296 6704 -3262
rect 6738 -3296 6764 -3262
rect 6678 -3330 6764 -3296
rect 6678 -3364 6704 -3330
rect 6738 -3364 6764 -3330
rect 6678 -3398 6764 -3364
rect 6678 -3432 6704 -3398
rect 6738 -3432 6764 -3398
rect 6678 -3466 6764 -3432
rect 6678 -3500 6704 -3466
rect 6738 -3500 6764 -3466
rect 6678 -3534 6764 -3500
rect 6678 -3568 6704 -3534
rect 6738 -3568 6764 -3534
rect 6678 -3602 6764 -3568
rect 6678 -3636 6704 -3602
rect 6738 -3636 6764 -3602
rect 6678 -3670 6764 -3636
rect 6678 -3704 6704 -3670
rect 6738 -3704 6764 -3670
rect 6678 -3738 6764 -3704
rect 6678 -3772 6704 -3738
rect 6738 -3772 6764 -3738
rect 6678 -3800 6764 -3772
rect 7872 -3460 7936 -3398
rect 7872 -3494 7898 -3460
rect 7932 -3494 7936 -3460
rect 7872 -3532 7936 -3494
rect 7872 -3566 7898 -3532
rect 7932 -3566 7936 -3532
rect 7872 -3600 7936 -3566
rect 7872 -3634 7898 -3600
rect 7932 -3634 7936 -3600
rect 7872 -3668 7936 -3634
rect 7872 -3702 7898 -3668
rect 7932 -3702 7936 -3668
rect 7872 -3736 7936 -3702
rect 7872 -3770 7898 -3736
rect 7932 -3770 7936 -3736
rect 7872 -3798 7936 -3770
rect 1968 -4440 2032 -4386
rect 1968 -4474 1994 -4440
rect 2028 -4474 2032 -4440
rect 1968 -4508 2032 -4474
rect 1968 -4542 1994 -4508
rect 2028 -4542 2032 -4508
rect 1968 -4576 2032 -4542
rect 1968 -4610 1994 -4576
rect 2028 -4610 2032 -4576
rect 1968 -4644 2032 -4610
rect 1968 -4678 1994 -4644
rect 2028 -4678 2032 -4644
rect 1968 -4712 2032 -4678
rect 1968 -4746 1994 -4712
rect 2028 -4746 2032 -4712
rect 1968 -4780 2032 -4746
rect 1968 -4814 1994 -4780
rect 2028 -4814 2032 -4780
rect 1968 -4848 2032 -4814
rect 1968 -4882 1994 -4848
rect 2028 -4882 2032 -4848
rect 1968 -4916 2032 -4882
rect 1968 -4950 1994 -4916
rect 2028 -4950 2032 -4916
rect 1968 -4984 2032 -4950
rect 1968 -5018 1994 -4984
rect 2028 -5018 2032 -4984
rect 1968 -5052 2032 -5018
rect 1968 -5086 1994 -5052
rect 2028 -5086 2032 -5052
rect 1968 -5120 2032 -5086
rect 1968 -5154 1994 -5120
rect 2028 -5154 2032 -5120
rect 1968 -5188 2032 -5154
rect 1968 -5222 1994 -5188
rect 2028 -5222 2032 -5188
rect 1968 -5256 2032 -5222
rect 1968 -5290 1994 -5256
rect 2028 -5290 2032 -5256
rect 1968 -5324 2032 -5290
rect 1968 -5358 1994 -5324
rect 2028 -5358 2032 -5324
rect 1968 -5386 2032 -5358
rect 2422 -4440 2508 -4386
rect 2422 -4474 2448 -4440
rect 2482 -4474 2508 -4440
rect 2422 -4508 2508 -4474
rect 2422 -4542 2448 -4508
rect 2482 -4542 2508 -4508
rect 2422 -4576 2508 -4542
rect 2422 -4610 2448 -4576
rect 2482 -4610 2508 -4576
rect 2422 -4644 2508 -4610
rect 2422 -4678 2448 -4644
rect 2482 -4678 2508 -4644
rect 2422 -4712 2508 -4678
rect 2422 -4746 2448 -4712
rect 2482 -4746 2508 -4712
rect 2422 -4780 2508 -4746
rect 2422 -4814 2448 -4780
rect 2482 -4814 2508 -4780
rect 2422 -4848 2508 -4814
rect 2422 -4882 2448 -4848
rect 2482 -4882 2508 -4848
rect 2422 -4916 2508 -4882
rect 2422 -4950 2448 -4916
rect 2482 -4950 2508 -4916
rect 2422 -4984 2508 -4950
rect 2422 -5018 2448 -4984
rect 2482 -5018 2508 -4984
rect 2422 -5052 2508 -5018
rect 2422 -5086 2448 -5052
rect 2482 -5086 2508 -5052
rect 2422 -5120 2508 -5086
rect 2422 -5154 2448 -5120
rect 2482 -5154 2508 -5120
rect 2422 -5188 2508 -5154
rect 2422 -5222 2448 -5188
rect 2482 -5222 2508 -5188
rect 2422 -5256 2508 -5222
rect 2422 -5290 2448 -5256
rect 2482 -5290 2508 -5256
rect 2422 -5324 2508 -5290
rect 2422 -5358 2448 -5324
rect 2482 -5358 2508 -5324
rect 2422 -5386 2508 -5358
rect 3486 -4440 3572 -4386
rect 3486 -4474 3512 -4440
rect 3546 -4474 3572 -4440
rect 3486 -4508 3572 -4474
rect 3486 -4542 3512 -4508
rect 3546 -4542 3572 -4508
rect 3486 -4576 3572 -4542
rect 3486 -4610 3512 -4576
rect 3546 -4610 3572 -4576
rect 3486 -4644 3572 -4610
rect 3486 -4678 3512 -4644
rect 3546 -4678 3572 -4644
rect 3486 -4712 3572 -4678
rect 3486 -4746 3512 -4712
rect 3546 -4746 3572 -4712
rect 3486 -4780 3572 -4746
rect 3486 -4814 3512 -4780
rect 3546 -4814 3572 -4780
rect 3486 -4848 3572 -4814
rect 3486 -4882 3512 -4848
rect 3546 -4882 3572 -4848
rect 3486 -4916 3572 -4882
rect 3486 -4950 3512 -4916
rect 3546 -4950 3572 -4916
rect 3486 -4984 3572 -4950
rect 3486 -5018 3512 -4984
rect 3546 -5018 3572 -4984
rect 3486 -5052 3572 -5018
rect 3486 -5086 3512 -5052
rect 3546 -5086 3572 -5052
rect 3486 -5120 3572 -5086
rect 3486 -5154 3512 -5120
rect 3546 -5154 3572 -5120
rect 3486 -5188 3572 -5154
rect 3486 -5222 3512 -5188
rect 3546 -5222 3572 -5188
rect 3486 -5256 3572 -5222
rect 3486 -5290 3512 -5256
rect 3546 -5290 3572 -5256
rect 3486 -5324 3572 -5290
rect 3486 -5358 3512 -5324
rect 3546 -5358 3572 -5324
rect 3486 -5386 3572 -5358
rect 4550 -4440 4636 -4386
rect 4550 -4474 4576 -4440
rect 4610 -4474 4636 -4440
rect 4550 -4508 4636 -4474
rect 4550 -4542 4576 -4508
rect 4610 -4542 4636 -4508
rect 4550 -4576 4636 -4542
rect 4550 -4610 4576 -4576
rect 4610 -4610 4636 -4576
rect 4550 -4644 4636 -4610
rect 4550 -4678 4576 -4644
rect 4610 -4678 4636 -4644
rect 4550 -4712 4636 -4678
rect 4550 -4746 4576 -4712
rect 4610 -4746 4636 -4712
rect 4550 -4780 4636 -4746
rect 4550 -4814 4576 -4780
rect 4610 -4814 4636 -4780
rect 4550 -4848 4636 -4814
rect 4550 -4882 4576 -4848
rect 4610 -4882 4636 -4848
rect 4550 -4916 4636 -4882
rect 4550 -4950 4576 -4916
rect 4610 -4950 4636 -4916
rect 4550 -4984 4636 -4950
rect 4550 -5018 4576 -4984
rect 4610 -5018 4636 -4984
rect 4550 -5052 4636 -5018
rect 4550 -5086 4576 -5052
rect 4610 -5086 4636 -5052
rect 4550 -5120 4636 -5086
rect 4550 -5154 4576 -5120
rect 4610 -5154 4636 -5120
rect 4550 -5188 4636 -5154
rect 4550 -5222 4576 -5188
rect 4610 -5222 4636 -5188
rect 4550 -5256 4636 -5222
rect 4550 -5290 4576 -5256
rect 4610 -5290 4636 -5256
rect 4550 -5324 4636 -5290
rect 4550 -5358 4576 -5324
rect 4610 -5358 4636 -5324
rect 4550 -5386 4636 -5358
rect 5614 -4440 5700 -4386
rect 5614 -4474 5640 -4440
rect 5674 -4474 5700 -4440
rect 5614 -4508 5700 -4474
rect 5614 -4542 5640 -4508
rect 5674 -4542 5700 -4508
rect 5614 -4576 5700 -4542
rect 5614 -4610 5640 -4576
rect 5674 -4610 5700 -4576
rect 5614 -4644 5700 -4610
rect 5614 -4678 5640 -4644
rect 5674 -4678 5700 -4644
rect 5614 -4712 5700 -4678
rect 5614 -4746 5640 -4712
rect 5674 -4746 5700 -4712
rect 5614 -4780 5700 -4746
rect 5614 -4814 5640 -4780
rect 5674 -4814 5700 -4780
rect 5614 -4848 5700 -4814
rect 5614 -4882 5640 -4848
rect 5674 -4882 5700 -4848
rect 5614 -4916 5700 -4882
rect 5614 -4950 5640 -4916
rect 5674 -4950 5700 -4916
rect 5614 -4984 5700 -4950
rect 5614 -5018 5640 -4984
rect 5674 -5018 5700 -4984
rect 5614 -5052 5700 -5018
rect 5614 -5086 5640 -5052
rect 5674 -5086 5700 -5052
rect 5614 -5120 5700 -5086
rect 5614 -5154 5640 -5120
rect 5674 -5154 5700 -5120
rect 5614 -5188 5700 -5154
rect 5614 -5222 5640 -5188
rect 5674 -5222 5700 -5188
rect 5614 -5256 5700 -5222
rect 5614 -5290 5640 -5256
rect 5674 -5290 5700 -5256
rect 5614 -5324 5700 -5290
rect 5614 -5358 5640 -5324
rect 5674 -5358 5700 -5324
rect 5614 -5386 5700 -5358
rect 6678 -4440 6764 -4386
rect 6678 -4474 6704 -4440
rect 6738 -4474 6764 -4440
rect 6678 -4508 6764 -4474
rect 6678 -4542 6704 -4508
rect 6738 -4542 6764 -4508
rect 6678 -4576 6764 -4542
rect 6678 -4610 6704 -4576
rect 6738 -4610 6764 -4576
rect 6678 -4644 6764 -4610
rect 6678 -4678 6704 -4644
rect 6738 -4678 6764 -4644
rect 6678 -4712 6764 -4678
rect 6678 -4746 6704 -4712
rect 6738 -4746 6764 -4712
rect 6678 -4780 6764 -4746
rect 6678 -4814 6704 -4780
rect 6738 -4814 6764 -4780
rect 6678 -4848 6764 -4814
rect 6678 -4882 6704 -4848
rect 6738 -4882 6764 -4848
rect 6678 -4916 6764 -4882
rect 6678 -4950 6704 -4916
rect 6738 -4950 6764 -4916
rect 6678 -4984 6764 -4950
rect 6678 -5018 6704 -4984
rect 6738 -5018 6764 -4984
rect 6678 -5052 6764 -5018
rect 6678 -5086 6704 -5052
rect 6738 -5086 6764 -5052
rect 6678 -5120 6764 -5086
rect 6678 -5154 6704 -5120
rect 6738 -5154 6764 -5120
rect 6678 -5188 6764 -5154
rect 6678 -5222 6704 -5188
rect 6738 -5222 6764 -5188
rect 6678 -5256 6764 -5222
rect 6678 -5290 6704 -5256
rect 6738 -5290 6764 -5256
rect 6678 -5324 6764 -5290
rect 6678 -5358 6704 -5324
rect 6738 -5358 6764 -5324
rect 6678 -5386 6764 -5358
rect 7872 -4448 7936 -4386
rect 7872 -4482 7898 -4448
rect 7932 -4482 7936 -4448
rect 7872 -4520 7936 -4482
rect 7872 -4554 7898 -4520
rect 7932 -4554 7936 -4520
rect 7872 -4588 7936 -4554
rect 7872 -4622 7898 -4588
rect 7932 -4622 7936 -4588
rect 7872 -4656 7936 -4622
rect 7872 -4690 7898 -4656
rect 7932 -4690 7936 -4656
rect 7872 -4724 7936 -4690
rect 7872 -4758 7898 -4724
rect 7932 -4758 7936 -4724
rect 7872 -4786 7936 -4758
rect 3796 -8868 3858 -8578
rect 4612 -8868 4674 -8578
rect 5428 -8868 5490 -8578
rect 6244 -8868 6306 -8578
rect 7060 -8868 7122 -8578
rect 3796 -9684 3858 -9394
rect 4612 -9684 4674 -9394
rect 5428 -9684 5490 -9394
rect 6244 -9684 6306 -9394
rect 7060 -9684 7122 -9394
<< psubdiffcont >>
rect 9584 -3336 9618 -3302
rect 9584 -3404 9618 -3370
rect 9584 -3472 9618 -3438
rect 9584 -3540 9618 -3506
rect 9584 -3608 9618 -3574
rect 9584 -3676 9618 -3642
rect 9584 -3744 9618 -3710
rect 9584 -3812 9618 -3778
rect 9584 -3880 9618 -3846
rect 9584 -3948 9618 -3914
rect 9584 -4016 9618 -3982
rect 9584 -4084 9618 -4050
rect 9584 -4152 9618 -4118
rect 9584 -4220 9618 -4186
rect 9584 -4492 9618 -4458
rect 9584 -4560 9618 -4526
rect 9584 -4628 9618 -4594
rect 9584 -4696 9618 -4662
rect 9584 -4764 9618 -4730
rect 9584 -4832 9618 -4798
rect 9584 -4900 9618 -4866
rect 9584 -4968 9618 -4934
rect 9584 -5036 9618 -5002
rect 9584 -5104 9618 -5070
rect 9584 -5172 9618 -5138
rect 9584 -5240 9618 -5206
rect 9584 -5308 9618 -5274
rect 9584 -5376 9618 -5342
rect 1642 -6234 1676 -6200
rect 1642 -6302 1676 -6268
rect 1642 -6370 1676 -6336
rect 1642 -6438 1676 -6404
rect 1642 -6506 1676 -6472
rect 1642 -6574 1676 -6540
rect 1642 -6642 1676 -6608
rect 1642 -6710 1676 -6676
rect 1642 -6778 1676 -6744
rect 1642 -6846 1676 -6812
rect 1642 -6914 1676 -6880
rect 1642 -6982 1676 -6948
rect 1642 -7050 1676 -7016
rect 1642 -7118 1676 -7084
rect 2706 -6234 2740 -6200
rect 2706 -6302 2740 -6268
rect 2706 -6370 2740 -6336
rect 2706 -6438 2740 -6404
rect 2706 -6506 2740 -6472
rect 2706 -6574 2740 -6540
rect 2706 -6642 2740 -6608
rect 2706 -6710 2740 -6676
rect 2706 -6778 2740 -6744
rect 2706 -6846 2740 -6812
rect 2706 -6914 2740 -6880
rect 2706 -6982 2740 -6948
rect 2706 -7050 2740 -7016
rect 2706 -7118 2740 -7084
rect 3770 -6234 3804 -6200
rect 3770 -6302 3804 -6268
rect 3770 -6370 3804 -6336
rect 3770 -6438 3804 -6404
rect 3770 -6506 3804 -6472
rect 3770 -6574 3804 -6540
rect 3770 -6642 3804 -6608
rect 3770 -6710 3804 -6676
rect 3770 -6778 3804 -6744
rect 3770 -6846 3804 -6812
rect 3770 -6914 3804 -6880
rect 3770 -6982 3804 -6948
rect 3770 -7050 3804 -7016
rect 3770 -7118 3804 -7084
rect 4834 -6234 4868 -6200
rect 4834 -6302 4868 -6268
rect 4834 -6370 4868 -6336
rect 4834 -6438 4868 -6404
rect 4834 -6506 4868 -6472
rect 4834 -6574 4868 -6540
rect 4834 -6642 4868 -6608
rect 4834 -6710 4868 -6676
rect 4834 -6778 4868 -6744
rect 4834 -6846 4868 -6812
rect 4834 -6914 4868 -6880
rect 4834 -6982 4868 -6948
rect 4834 -7050 4868 -7016
rect 4834 -7118 4868 -7084
rect 5994 -6234 6028 -6200
rect 5994 -6302 6028 -6268
rect 5994 -6370 6028 -6336
rect 5994 -6438 6028 -6404
rect 5994 -6506 6028 -6472
rect 5994 -6574 6028 -6540
rect 5994 -6642 6028 -6608
rect 5994 -6710 6028 -6676
rect 5994 -6778 6028 -6744
rect 5994 -6846 6028 -6812
rect 5994 -6914 6028 -6880
rect 5994 -6982 6028 -6948
rect 5994 -7050 6028 -7016
rect 5994 -7118 6028 -7084
rect 7058 -6234 7092 -6200
rect 7058 -6302 7092 -6268
rect 7058 -6370 7092 -6336
rect 7058 -6438 7092 -6404
rect 7058 -6506 7092 -6472
rect 7058 -6574 7092 -6540
rect 7058 -6642 7092 -6608
rect 7058 -6710 7092 -6676
rect 7058 -6778 7092 -6744
rect 7058 -6846 7092 -6812
rect 7058 -6914 7092 -6880
rect 7058 -6982 7092 -6948
rect 7058 -7050 7092 -7016
rect 7058 -7118 7092 -7084
rect 8122 -6234 8156 -6200
rect 8122 -6302 8156 -6268
rect 8122 -6370 8156 -6336
rect 8122 -6438 8156 -6404
rect 8122 -6506 8156 -6472
rect 8122 -6574 8156 -6540
rect 8122 -6642 8156 -6608
rect 8122 -6710 8156 -6676
rect 8122 -6778 8156 -6744
rect 8122 -6846 8156 -6812
rect 8122 -6914 8156 -6880
rect 8122 -6982 8156 -6948
rect 8122 -7050 8156 -7016
rect 8122 -7118 8156 -7084
rect 8962 -6150 9042 -5978
rect 8962 -6494 9042 -6322
rect 8962 -6838 9042 -6666
rect 8962 -7182 9042 -7010
rect 1170 -7590 1250 -7418
rect 1170 -7934 1250 -7762
rect 8962 -7526 9042 -7354
rect 8962 -7870 9042 -7698
rect 1170 -8278 1250 -8106
<< nsubdiffcont >>
rect 1994 -2888 2028 -2854
rect 1994 -2956 2028 -2922
rect 1994 -3024 2028 -2990
rect 1994 -3092 2028 -3058
rect 1994 -3160 2028 -3126
rect 1994 -3228 2028 -3194
rect 1994 -3296 2028 -3262
rect 1994 -3364 2028 -3330
rect 1994 -3432 2028 -3398
rect 1994 -3500 2028 -3466
rect 1994 -3568 2028 -3534
rect 1994 -3636 2028 -3602
rect 1994 -3704 2028 -3670
rect 1994 -3772 2028 -3738
rect 2448 -2888 2482 -2854
rect 2448 -2956 2482 -2922
rect 2448 -3024 2482 -2990
rect 2448 -3092 2482 -3058
rect 2448 -3160 2482 -3126
rect 2448 -3228 2482 -3194
rect 2448 -3296 2482 -3262
rect 2448 -3364 2482 -3330
rect 2448 -3432 2482 -3398
rect 2448 -3500 2482 -3466
rect 2448 -3568 2482 -3534
rect 2448 -3636 2482 -3602
rect 2448 -3704 2482 -3670
rect 2448 -3772 2482 -3738
rect 3512 -2888 3546 -2854
rect 3512 -2956 3546 -2922
rect 3512 -3024 3546 -2990
rect 3512 -3092 3546 -3058
rect 3512 -3160 3546 -3126
rect 3512 -3228 3546 -3194
rect 3512 -3296 3546 -3262
rect 3512 -3364 3546 -3330
rect 3512 -3432 3546 -3398
rect 3512 -3500 3546 -3466
rect 3512 -3568 3546 -3534
rect 3512 -3636 3546 -3602
rect 3512 -3704 3546 -3670
rect 3512 -3772 3546 -3738
rect 4576 -2888 4610 -2854
rect 4576 -2956 4610 -2922
rect 4576 -3024 4610 -2990
rect 4576 -3092 4610 -3058
rect 4576 -3160 4610 -3126
rect 4576 -3228 4610 -3194
rect 4576 -3296 4610 -3262
rect 4576 -3364 4610 -3330
rect 4576 -3432 4610 -3398
rect 4576 -3500 4610 -3466
rect 4576 -3568 4610 -3534
rect 4576 -3636 4610 -3602
rect 4576 -3704 4610 -3670
rect 4576 -3772 4610 -3738
rect 5640 -2888 5674 -2854
rect 5640 -2956 5674 -2922
rect 5640 -3024 5674 -2990
rect 5640 -3092 5674 -3058
rect 5640 -3160 5674 -3126
rect 5640 -3228 5674 -3194
rect 5640 -3296 5674 -3262
rect 5640 -3364 5674 -3330
rect 5640 -3432 5674 -3398
rect 5640 -3500 5674 -3466
rect 5640 -3568 5674 -3534
rect 5640 -3636 5674 -3602
rect 5640 -3704 5674 -3670
rect 5640 -3772 5674 -3738
rect 6704 -2888 6738 -2854
rect 6704 -2956 6738 -2922
rect 6704 -3024 6738 -2990
rect 6704 -3092 6738 -3058
rect 6704 -3160 6738 -3126
rect 6704 -3228 6738 -3194
rect 6704 -3296 6738 -3262
rect 6704 -3364 6738 -3330
rect 6704 -3432 6738 -3398
rect 6704 -3500 6738 -3466
rect 6704 -3568 6738 -3534
rect 6704 -3636 6738 -3602
rect 6704 -3704 6738 -3670
rect 6704 -3772 6738 -3738
rect 7898 -3494 7932 -3460
rect 7898 -3566 7932 -3532
rect 7898 -3634 7932 -3600
rect 7898 -3702 7932 -3668
rect 7898 -3770 7932 -3736
rect 1994 -4474 2028 -4440
rect 1994 -4542 2028 -4508
rect 1994 -4610 2028 -4576
rect 1994 -4678 2028 -4644
rect 1994 -4746 2028 -4712
rect 1994 -4814 2028 -4780
rect 1994 -4882 2028 -4848
rect 1994 -4950 2028 -4916
rect 1994 -5018 2028 -4984
rect 1994 -5086 2028 -5052
rect 1994 -5154 2028 -5120
rect 1994 -5222 2028 -5188
rect 1994 -5290 2028 -5256
rect 1994 -5358 2028 -5324
rect 2448 -4474 2482 -4440
rect 2448 -4542 2482 -4508
rect 2448 -4610 2482 -4576
rect 2448 -4678 2482 -4644
rect 2448 -4746 2482 -4712
rect 2448 -4814 2482 -4780
rect 2448 -4882 2482 -4848
rect 2448 -4950 2482 -4916
rect 2448 -5018 2482 -4984
rect 2448 -5086 2482 -5052
rect 2448 -5154 2482 -5120
rect 2448 -5222 2482 -5188
rect 2448 -5290 2482 -5256
rect 2448 -5358 2482 -5324
rect 3512 -4474 3546 -4440
rect 3512 -4542 3546 -4508
rect 3512 -4610 3546 -4576
rect 3512 -4678 3546 -4644
rect 3512 -4746 3546 -4712
rect 3512 -4814 3546 -4780
rect 3512 -4882 3546 -4848
rect 3512 -4950 3546 -4916
rect 3512 -5018 3546 -4984
rect 3512 -5086 3546 -5052
rect 3512 -5154 3546 -5120
rect 3512 -5222 3546 -5188
rect 3512 -5290 3546 -5256
rect 3512 -5358 3546 -5324
rect 4576 -4474 4610 -4440
rect 4576 -4542 4610 -4508
rect 4576 -4610 4610 -4576
rect 4576 -4678 4610 -4644
rect 4576 -4746 4610 -4712
rect 4576 -4814 4610 -4780
rect 4576 -4882 4610 -4848
rect 4576 -4950 4610 -4916
rect 4576 -5018 4610 -4984
rect 4576 -5086 4610 -5052
rect 4576 -5154 4610 -5120
rect 4576 -5222 4610 -5188
rect 4576 -5290 4610 -5256
rect 4576 -5358 4610 -5324
rect 5640 -4474 5674 -4440
rect 5640 -4542 5674 -4508
rect 5640 -4610 5674 -4576
rect 5640 -4678 5674 -4644
rect 5640 -4746 5674 -4712
rect 5640 -4814 5674 -4780
rect 5640 -4882 5674 -4848
rect 5640 -4950 5674 -4916
rect 5640 -5018 5674 -4984
rect 5640 -5086 5674 -5052
rect 5640 -5154 5674 -5120
rect 5640 -5222 5674 -5188
rect 5640 -5290 5674 -5256
rect 5640 -5358 5674 -5324
rect 6704 -4474 6738 -4440
rect 6704 -4542 6738 -4508
rect 6704 -4610 6738 -4576
rect 6704 -4678 6738 -4644
rect 6704 -4746 6738 -4712
rect 6704 -4814 6738 -4780
rect 6704 -4882 6738 -4848
rect 6704 -4950 6738 -4916
rect 6704 -5018 6738 -4984
rect 6704 -5086 6738 -5052
rect 6704 -5154 6738 -5120
rect 6704 -5222 6738 -5188
rect 6704 -5290 6738 -5256
rect 6704 -5358 6738 -5324
rect 7898 -4482 7932 -4448
rect 7898 -4554 7932 -4520
rect 7898 -4622 7932 -4588
rect 7898 -4690 7932 -4656
rect 7898 -4758 7932 -4724
<< locali >>
rect 1994 -2812 2028 -2796
rect 1994 -3804 2028 -3788
rect 2448 -2812 2482 -2796
rect 2448 -3804 2482 -3788
rect 3512 -2812 3546 -2796
rect 3512 -3804 3546 -3788
rect 4576 -2812 4610 -2796
rect 4576 -3804 4610 -3788
rect 5640 -2812 5674 -2796
rect 5640 -3804 5674 -3788
rect 6704 -2812 6738 -2796
rect 9584 -3260 9618 -3244
rect 6704 -3804 6738 -3788
rect 7898 -3410 7932 -3394
rect 7898 -3802 7932 -3786
rect 9584 -4252 9618 -4236
rect 1994 -4398 2028 -4382
rect 1994 -5390 2028 -5374
rect 2448 -4398 2482 -4382
rect 2448 -5390 2482 -5374
rect 3512 -4398 3546 -4382
rect 3512 -5386 3546 -5374
rect 4576 -4398 4610 -4382
rect 4576 -5386 4610 -5374
rect 5640 -4398 5674 -4382
rect 5640 -5386 5674 -5374
rect 6704 -4398 6738 -4382
rect 7898 -4398 7932 -4382
rect 7898 -4786 7932 -4774
rect 9584 -4416 9618 -4400
rect 6704 -5386 6738 -5374
rect 9584 -5408 9618 -5392
rect 8962 -5978 9042 -5886
rect 1642 -6200 1676 -6142
rect 1642 -6268 1676 -6234
rect 1642 -6336 1676 -6302
rect 1642 -6404 1676 -6370
rect 1642 -6472 1676 -6438
rect 1642 -6540 1676 -6506
rect 1642 -6608 1676 -6574
rect 1642 -6676 1676 -6642
rect 1642 -6744 1676 -6710
rect 1642 -6812 1676 -6778
rect 1642 -6880 1676 -6846
rect 1642 -6948 1676 -6914
rect 1642 -7016 1676 -6982
rect 1642 -7084 1676 -7050
rect 1642 -7150 1676 -7118
rect 2706 -6200 2740 -6142
rect 2706 -6268 2740 -6234
rect 2706 -6336 2740 -6302
rect 2706 -6404 2740 -6370
rect 2706 -6472 2740 -6438
rect 2706 -6540 2740 -6506
rect 2706 -6608 2740 -6574
rect 2706 -6676 2740 -6642
rect 2706 -6744 2740 -6710
rect 2706 -6812 2740 -6778
rect 2706 -6880 2740 -6846
rect 2706 -6948 2740 -6914
rect 2706 -7016 2740 -6982
rect 2706 -7084 2740 -7050
rect 2706 -7150 2740 -7118
rect 3770 -6200 3804 -6142
rect 3770 -6268 3804 -6234
rect 3770 -6336 3804 -6302
rect 3770 -6404 3804 -6370
rect 3770 -6472 3804 -6438
rect 3770 -6540 3804 -6506
rect 3770 -6608 3804 -6574
rect 3770 -6676 3804 -6642
rect 3770 -6744 3804 -6710
rect 3770 -6812 3804 -6778
rect 3770 -6880 3804 -6846
rect 3770 -6948 3804 -6914
rect 3770 -7016 3804 -6982
rect 3770 -7084 3804 -7050
rect 3770 -7150 3804 -7118
rect 4834 -6200 4868 -6142
rect 4834 -6268 4868 -6234
rect 4834 -6336 4868 -6302
rect 4834 -6404 4868 -6370
rect 4834 -6472 4868 -6438
rect 4834 -6540 4868 -6506
rect 4834 -6608 4868 -6574
rect 4834 -6676 4868 -6642
rect 4834 -6744 4868 -6710
rect 4834 -6812 4868 -6778
rect 4834 -6880 4868 -6846
rect 4834 -6948 4868 -6914
rect 4834 -7016 4868 -6982
rect 4834 -7084 4868 -7050
rect 4834 -7150 4868 -7118
rect 5994 -6158 6028 -6142
rect 5994 -7150 6028 -7134
rect 7058 -6158 7092 -6142
rect 7058 -7150 7092 -7134
rect 8122 -6158 8156 -6142
rect 8122 -7150 8156 -7134
rect 1170 -7418 1250 -7260
rect 8962 -7950 9042 -7870
rect 1170 -8312 1250 -8278
<< viali >>
rect 1994 -2854 2028 -2812
rect 1994 -2888 2028 -2854
rect 1994 -2922 2028 -2888
rect 1994 -2956 2028 -2922
rect 1994 -2990 2028 -2956
rect 1994 -3024 2028 -2990
rect 1994 -3058 2028 -3024
rect 1994 -3092 2028 -3058
rect 1994 -3126 2028 -3092
rect 1994 -3160 2028 -3126
rect 1994 -3194 2028 -3160
rect 1994 -3228 2028 -3194
rect 1994 -3262 2028 -3228
rect 1994 -3296 2028 -3262
rect 1994 -3330 2028 -3296
rect 1994 -3364 2028 -3330
rect 1994 -3398 2028 -3364
rect 1994 -3432 2028 -3398
rect 1994 -3466 2028 -3432
rect 1994 -3500 2028 -3466
rect 1994 -3534 2028 -3500
rect 1994 -3568 2028 -3534
rect 1994 -3602 2028 -3568
rect 1994 -3636 2028 -3602
rect 1994 -3670 2028 -3636
rect 1994 -3704 2028 -3670
rect 1994 -3738 2028 -3704
rect 1994 -3772 2028 -3738
rect 1994 -3788 2028 -3772
rect 2448 -2854 2482 -2812
rect 2448 -2888 2482 -2854
rect 2448 -2922 2482 -2888
rect 2448 -2956 2482 -2922
rect 2448 -2990 2482 -2956
rect 2448 -3024 2482 -2990
rect 2448 -3058 2482 -3024
rect 2448 -3092 2482 -3058
rect 2448 -3126 2482 -3092
rect 2448 -3160 2482 -3126
rect 2448 -3194 2482 -3160
rect 2448 -3228 2482 -3194
rect 2448 -3262 2482 -3228
rect 2448 -3296 2482 -3262
rect 2448 -3330 2482 -3296
rect 2448 -3364 2482 -3330
rect 2448 -3398 2482 -3364
rect 2448 -3432 2482 -3398
rect 2448 -3466 2482 -3432
rect 2448 -3500 2482 -3466
rect 2448 -3534 2482 -3500
rect 2448 -3568 2482 -3534
rect 2448 -3602 2482 -3568
rect 2448 -3636 2482 -3602
rect 2448 -3670 2482 -3636
rect 2448 -3704 2482 -3670
rect 2448 -3738 2482 -3704
rect 2448 -3772 2482 -3738
rect 2448 -3788 2482 -3772
rect 3512 -2854 3546 -2812
rect 3512 -2888 3546 -2854
rect 3512 -2922 3546 -2888
rect 3512 -2956 3546 -2922
rect 3512 -2990 3546 -2956
rect 3512 -3024 3546 -2990
rect 3512 -3058 3546 -3024
rect 3512 -3092 3546 -3058
rect 3512 -3126 3546 -3092
rect 3512 -3160 3546 -3126
rect 3512 -3194 3546 -3160
rect 3512 -3228 3546 -3194
rect 3512 -3262 3546 -3228
rect 3512 -3296 3546 -3262
rect 3512 -3330 3546 -3296
rect 3512 -3364 3546 -3330
rect 3512 -3398 3546 -3364
rect 3512 -3432 3546 -3398
rect 3512 -3466 3546 -3432
rect 3512 -3500 3546 -3466
rect 3512 -3534 3546 -3500
rect 3512 -3568 3546 -3534
rect 3512 -3602 3546 -3568
rect 3512 -3636 3546 -3602
rect 3512 -3670 3546 -3636
rect 3512 -3704 3546 -3670
rect 3512 -3738 3546 -3704
rect 3512 -3772 3546 -3738
rect 3512 -3788 3546 -3772
rect 4576 -2854 4610 -2812
rect 4576 -2888 4610 -2854
rect 4576 -2922 4610 -2888
rect 4576 -2956 4610 -2922
rect 4576 -2990 4610 -2956
rect 4576 -3024 4610 -2990
rect 4576 -3058 4610 -3024
rect 4576 -3092 4610 -3058
rect 4576 -3126 4610 -3092
rect 4576 -3160 4610 -3126
rect 4576 -3194 4610 -3160
rect 4576 -3228 4610 -3194
rect 4576 -3262 4610 -3228
rect 4576 -3296 4610 -3262
rect 4576 -3330 4610 -3296
rect 4576 -3364 4610 -3330
rect 4576 -3398 4610 -3364
rect 4576 -3432 4610 -3398
rect 4576 -3466 4610 -3432
rect 4576 -3500 4610 -3466
rect 4576 -3534 4610 -3500
rect 4576 -3568 4610 -3534
rect 4576 -3602 4610 -3568
rect 4576 -3636 4610 -3602
rect 4576 -3670 4610 -3636
rect 4576 -3704 4610 -3670
rect 4576 -3738 4610 -3704
rect 4576 -3772 4610 -3738
rect 4576 -3788 4610 -3772
rect 5640 -2854 5674 -2812
rect 5640 -2888 5674 -2854
rect 5640 -2922 5674 -2888
rect 5640 -2956 5674 -2922
rect 5640 -2990 5674 -2956
rect 5640 -3024 5674 -2990
rect 5640 -3058 5674 -3024
rect 5640 -3092 5674 -3058
rect 5640 -3126 5674 -3092
rect 5640 -3160 5674 -3126
rect 5640 -3194 5674 -3160
rect 5640 -3228 5674 -3194
rect 5640 -3262 5674 -3228
rect 5640 -3296 5674 -3262
rect 5640 -3330 5674 -3296
rect 5640 -3364 5674 -3330
rect 5640 -3398 5674 -3364
rect 5640 -3432 5674 -3398
rect 5640 -3466 5674 -3432
rect 5640 -3500 5674 -3466
rect 5640 -3534 5674 -3500
rect 5640 -3568 5674 -3534
rect 5640 -3602 5674 -3568
rect 5640 -3636 5674 -3602
rect 5640 -3670 5674 -3636
rect 5640 -3704 5674 -3670
rect 5640 -3738 5674 -3704
rect 5640 -3772 5674 -3738
rect 5640 -3788 5674 -3772
rect 6704 -2854 6738 -2812
rect 6704 -2888 6738 -2854
rect 6704 -2922 6738 -2888
rect 6704 -2956 6738 -2922
rect 6704 -2990 6738 -2956
rect 6704 -3024 6738 -2990
rect 6704 -3058 6738 -3024
rect 6704 -3092 6738 -3058
rect 6704 -3126 6738 -3092
rect 6704 -3160 6738 -3126
rect 6704 -3194 6738 -3160
rect 6704 -3228 6738 -3194
rect 6704 -3262 6738 -3228
rect 6704 -3296 6738 -3262
rect 6704 -3330 6738 -3296
rect 6704 -3364 6738 -3330
rect 6704 -3398 6738 -3364
rect 9584 -3302 9618 -3260
rect 9584 -3336 9618 -3302
rect 9584 -3370 9618 -3336
rect 6704 -3432 6738 -3398
rect 6704 -3466 6738 -3432
rect 6704 -3500 6738 -3466
rect 6704 -3534 6738 -3500
rect 6704 -3568 6738 -3534
rect 6704 -3602 6738 -3568
rect 6704 -3636 6738 -3602
rect 6704 -3670 6738 -3636
rect 6704 -3704 6738 -3670
rect 6704 -3738 6738 -3704
rect 6704 -3772 6738 -3738
rect 6704 -3788 6738 -3772
rect 7898 -3460 7932 -3410
rect 7898 -3494 7932 -3460
rect 7898 -3532 7932 -3494
rect 7898 -3566 7932 -3532
rect 7898 -3600 7932 -3566
rect 7898 -3634 7932 -3600
rect 7898 -3668 7932 -3634
rect 7898 -3702 7932 -3668
rect 7898 -3736 7932 -3702
rect 7898 -3770 7932 -3736
rect 7898 -3786 7932 -3770
rect 9584 -3404 9618 -3370
rect 9584 -3438 9618 -3404
rect 9584 -3472 9618 -3438
rect 9584 -3506 9618 -3472
rect 9584 -3540 9618 -3506
rect 9584 -3574 9618 -3540
rect 9584 -3608 9618 -3574
rect 9584 -3642 9618 -3608
rect 9584 -3676 9618 -3642
rect 9584 -3710 9618 -3676
rect 9584 -3744 9618 -3710
rect 9584 -3778 9618 -3744
rect 9584 -3812 9618 -3778
rect 9584 -3846 9618 -3812
rect 9584 -3880 9618 -3846
rect 9584 -3914 9618 -3880
rect 9584 -3948 9618 -3914
rect 9584 -3982 9618 -3948
rect 9584 -4016 9618 -3982
rect 9584 -4050 9618 -4016
rect 9584 -4084 9618 -4050
rect 9584 -4118 9618 -4084
rect 9584 -4152 9618 -4118
rect 9584 -4186 9618 -4152
rect 9584 -4220 9618 -4186
rect 9584 -4236 9618 -4220
rect 1994 -4440 2028 -4398
rect 1994 -4474 2028 -4440
rect 1994 -4508 2028 -4474
rect 1994 -4542 2028 -4508
rect 1994 -4576 2028 -4542
rect 1994 -4610 2028 -4576
rect 1994 -4644 2028 -4610
rect 1994 -4678 2028 -4644
rect 1994 -4712 2028 -4678
rect 1994 -4746 2028 -4712
rect 1994 -4780 2028 -4746
rect 1994 -4814 2028 -4780
rect 1994 -4848 2028 -4814
rect 1994 -4882 2028 -4848
rect 1994 -4916 2028 -4882
rect 1994 -4950 2028 -4916
rect 1994 -4984 2028 -4950
rect 1994 -5018 2028 -4984
rect 1994 -5052 2028 -5018
rect 1994 -5086 2028 -5052
rect 1994 -5120 2028 -5086
rect 1994 -5154 2028 -5120
rect 1994 -5188 2028 -5154
rect 1994 -5222 2028 -5188
rect 1994 -5256 2028 -5222
rect 1994 -5290 2028 -5256
rect 1994 -5324 2028 -5290
rect 1994 -5358 2028 -5324
rect 1994 -5374 2028 -5358
rect 2448 -4440 2482 -4398
rect 2448 -4474 2482 -4440
rect 2448 -4508 2482 -4474
rect 2448 -4542 2482 -4508
rect 2448 -4576 2482 -4542
rect 2448 -4610 2482 -4576
rect 2448 -4644 2482 -4610
rect 2448 -4678 2482 -4644
rect 2448 -4712 2482 -4678
rect 2448 -4746 2482 -4712
rect 2448 -4780 2482 -4746
rect 2448 -4814 2482 -4780
rect 2448 -4848 2482 -4814
rect 2448 -4882 2482 -4848
rect 2448 -4916 2482 -4882
rect 2448 -4950 2482 -4916
rect 2448 -4984 2482 -4950
rect 2448 -5018 2482 -4984
rect 2448 -5052 2482 -5018
rect 2448 -5086 2482 -5052
rect 2448 -5120 2482 -5086
rect 2448 -5154 2482 -5120
rect 2448 -5188 2482 -5154
rect 2448 -5222 2482 -5188
rect 2448 -5256 2482 -5222
rect 2448 -5290 2482 -5256
rect 2448 -5324 2482 -5290
rect 2448 -5358 2482 -5324
rect 2448 -5374 2482 -5358
rect 3512 -4440 3546 -4398
rect 3512 -4474 3546 -4440
rect 3512 -4508 3546 -4474
rect 3512 -4542 3546 -4508
rect 3512 -4576 3546 -4542
rect 3512 -4610 3546 -4576
rect 3512 -4644 3546 -4610
rect 3512 -4678 3546 -4644
rect 3512 -4712 3546 -4678
rect 3512 -4746 3546 -4712
rect 3512 -4780 3546 -4746
rect 3512 -4814 3546 -4780
rect 3512 -4848 3546 -4814
rect 3512 -4882 3546 -4848
rect 3512 -4916 3546 -4882
rect 3512 -4950 3546 -4916
rect 3512 -4984 3546 -4950
rect 3512 -5018 3546 -4984
rect 3512 -5052 3546 -5018
rect 3512 -5086 3546 -5052
rect 3512 -5120 3546 -5086
rect 3512 -5154 3546 -5120
rect 3512 -5188 3546 -5154
rect 3512 -5222 3546 -5188
rect 3512 -5256 3546 -5222
rect 3512 -5290 3546 -5256
rect 3512 -5324 3546 -5290
rect 3512 -5358 3546 -5324
rect 3512 -5374 3546 -5358
rect 4576 -4440 4610 -4398
rect 4576 -4474 4610 -4440
rect 4576 -4508 4610 -4474
rect 4576 -4542 4610 -4508
rect 4576 -4576 4610 -4542
rect 4576 -4610 4610 -4576
rect 4576 -4644 4610 -4610
rect 4576 -4678 4610 -4644
rect 4576 -4712 4610 -4678
rect 4576 -4746 4610 -4712
rect 4576 -4780 4610 -4746
rect 4576 -4814 4610 -4780
rect 4576 -4848 4610 -4814
rect 4576 -4882 4610 -4848
rect 4576 -4916 4610 -4882
rect 4576 -4950 4610 -4916
rect 4576 -4984 4610 -4950
rect 4576 -5018 4610 -4984
rect 4576 -5052 4610 -5018
rect 4576 -5086 4610 -5052
rect 4576 -5120 4610 -5086
rect 4576 -5154 4610 -5120
rect 4576 -5188 4610 -5154
rect 4576 -5222 4610 -5188
rect 4576 -5256 4610 -5222
rect 4576 -5290 4610 -5256
rect 4576 -5324 4610 -5290
rect 4576 -5358 4610 -5324
rect 4576 -5374 4610 -5358
rect 5640 -4440 5674 -4398
rect 5640 -4474 5674 -4440
rect 5640 -4508 5674 -4474
rect 5640 -4542 5674 -4508
rect 5640 -4576 5674 -4542
rect 5640 -4610 5674 -4576
rect 5640 -4644 5674 -4610
rect 5640 -4678 5674 -4644
rect 5640 -4712 5674 -4678
rect 5640 -4746 5674 -4712
rect 5640 -4780 5674 -4746
rect 5640 -4814 5674 -4780
rect 5640 -4848 5674 -4814
rect 5640 -4882 5674 -4848
rect 5640 -4916 5674 -4882
rect 5640 -4950 5674 -4916
rect 5640 -4984 5674 -4950
rect 5640 -5018 5674 -4984
rect 5640 -5052 5674 -5018
rect 5640 -5086 5674 -5052
rect 5640 -5120 5674 -5086
rect 5640 -5154 5674 -5120
rect 5640 -5188 5674 -5154
rect 5640 -5222 5674 -5188
rect 5640 -5256 5674 -5222
rect 5640 -5290 5674 -5256
rect 5640 -5324 5674 -5290
rect 5640 -5358 5674 -5324
rect 5640 -5374 5674 -5358
rect 6704 -4440 6738 -4398
rect 6704 -4474 6738 -4440
rect 6704 -4508 6738 -4474
rect 6704 -4542 6738 -4508
rect 6704 -4576 6738 -4542
rect 6704 -4610 6738 -4576
rect 6704 -4644 6738 -4610
rect 6704 -4678 6738 -4644
rect 6704 -4712 6738 -4678
rect 6704 -4746 6738 -4712
rect 6704 -4780 6738 -4746
rect 6704 -4814 6738 -4780
rect 7898 -4448 7932 -4398
rect 7898 -4482 7932 -4448
rect 7898 -4520 7932 -4482
rect 7898 -4554 7932 -4520
rect 7898 -4588 7932 -4554
rect 7898 -4622 7932 -4588
rect 7898 -4656 7932 -4622
rect 7898 -4690 7932 -4656
rect 7898 -4724 7932 -4690
rect 7898 -4758 7932 -4724
rect 7898 -4774 7932 -4758
rect 9584 -4458 9618 -4416
rect 9584 -4492 9618 -4458
rect 9584 -4526 9618 -4492
rect 9584 -4560 9618 -4526
rect 9584 -4594 9618 -4560
rect 9584 -4628 9618 -4594
rect 9584 -4662 9618 -4628
rect 9584 -4696 9618 -4662
rect 9584 -4730 9618 -4696
rect 9584 -4764 9618 -4730
rect 6704 -4848 6738 -4814
rect 6704 -4882 6738 -4848
rect 6704 -4916 6738 -4882
rect 6704 -4950 6738 -4916
rect 6704 -4984 6738 -4950
rect 6704 -5018 6738 -4984
rect 6704 -5052 6738 -5018
rect 6704 -5086 6738 -5052
rect 6704 -5120 6738 -5086
rect 6704 -5154 6738 -5120
rect 6704 -5188 6738 -5154
rect 6704 -5222 6738 -5188
rect 6704 -5256 6738 -5222
rect 6704 -5290 6738 -5256
rect 6704 -5324 6738 -5290
rect 6704 -5358 6738 -5324
rect 6704 -5374 6738 -5358
rect 9584 -4798 9618 -4764
rect 9584 -4832 9618 -4798
rect 9584 -4866 9618 -4832
rect 9584 -4900 9618 -4866
rect 9584 -4934 9618 -4900
rect 9584 -4968 9618 -4934
rect 9584 -5002 9618 -4968
rect 9584 -5036 9618 -5002
rect 9584 -5070 9618 -5036
rect 9584 -5104 9618 -5070
rect 9584 -5138 9618 -5104
rect 9584 -5172 9618 -5138
rect 9584 -5206 9618 -5172
rect 9584 -5240 9618 -5206
rect 9584 -5274 9618 -5240
rect 9584 -5308 9618 -5274
rect 9584 -5342 9618 -5308
rect 9584 -5376 9618 -5342
rect 9584 -5392 9618 -5376
rect 5994 -6200 6028 -6158
rect 5994 -6234 6028 -6200
rect 5994 -6268 6028 -6234
rect 5994 -6302 6028 -6268
rect 5994 -6336 6028 -6302
rect 5994 -6370 6028 -6336
rect 5994 -6404 6028 -6370
rect 5994 -6438 6028 -6404
rect 5994 -6472 6028 -6438
rect 5994 -6506 6028 -6472
rect 5994 -6540 6028 -6506
rect 5994 -6574 6028 -6540
rect 5994 -6608 6028 -6574
rect 5994 -6642 6028 -6608
rect 5994 -6676 6028 -6642
rect 5994 -6710 6028 -6676
rect 5994 -6744 6028 -6710
rect 5994 -6778 6028 -6744
rect 5994 -6812 6028 -6778
rect 5994 -6846 6028 -6812
rect 5994 -6880 6028 -6846
rect 5994 -6914 6028 -6880
rect 5994 -6948 6028 -6914
rect 5994 -6982 6028 -6948
rect 5994 -7016 6028 -6982
rect 5994 -7050 6028 -7016
rect 5994 -7084 6028 -7050
rect 5994 -7118 6028 -7084
rect 5994 -7134 6028 -7118
rect 7058 -6200 7092 -6158
rect 7058 -6234 7092 -6200
rect 7058 -6268 7092 -6234
rect 7058 -6302 7092 -6268
rect 7058 -6336 7092 -6302
rect 7058 -6370 7092 -6336
rect 7058 -6404 7092 -6370
rect 7058 -6438 7092 -6404
rect 7058 -6472 7092 -6438
rect 7058 -6506 7092 -6472
rect 7058 -6540 7092 -6506
rect 7058 -6574 7092 -6540
rect 7058 -6608 7092 -6574
rect 7058 -6642 7092 -6608
rect 7058 -6676 7092 -6642
rect 7058 -6710 7092 -6676
rect 7058 -6744 7092 -6710
rect 7058 -6778 7092 -6744
rect 7058 -6812 7092 -6778
rect 7058 -6846 7092 -6812
rect 7058 -6880 7092 -6846
rect 7058 -6914 7092 -6880
rect 7058 -6948 7092 -6914
rect 7058 -6982 7092 -6948
rect 7058 -7016 7092 -6982
rect 7058 -7050 7092 -7016
rect 7058 -7084 7092 -7050
rect 7058 -7118 7092 -7084
rect 7058 -7134 7092 -7118
rect 8122 -6200 8156 -6158
rect 8122 -6234 8156 -6200
rect 8122 -6268 8156 -6234
rect 8122 -6302 8156 -6268
rect 8122 -6336 8156 -6302
rect 8122 -6370 8156 -6336
rect 8122 -6404 8156 -6370
rect 8122 -6438 8156 -6404
rect 8122 -6472 8156 -6438
rect 8122 -6506 8156 -6472
rect 8122 -6540 8156 -6506
rect 8122 -6574 8156 -6540
rect 8122 -6608 8156 -6574
rect 8122 -6642 8156 -6608
rect 8122 -6676 8156 -6642
rect 8122 -6710 8156 -6676
rect 8122 -6744 8156 -6710
rect 8122 -6778 8156 -6744
rect 8122 -6812 8156 -6778
rect 8122 -6846 8156 -6812
rect 8122 -6880 8156 -6846
rect 8122 -6914 8156 -6880
rect 8122 -6948 8156 -6914
rect 8122 -6982 8156 -6948
rect 8122 -7016 8156 -6982
rect 8122 -7050 8156 -7016
rect 8122 -7084 8156 -7050
rect 8122 -7118 8156 -7084
rect 8122 -7134 8156 -7118
rect 8962 -6150 9042 -5978
rect 8962 -6322 9042 -6150
rect 8962 -6494 9042 -6322
rect 8962 -6666 9042 -6494
rect 8962 -6838 9042 -6666
rect 8962 -7010 9042 -6838
rect 8962 -7182 9042 -7010
rect 1170 -7590 1250 -7418
rect 1170 -7762 1250 -7590
rect 1170 -7934 1250 -7762
rect 1170 -8106 1250 -7934
rect 8962 -7354 9042 -7182
rect 8962 -7526 9042 -7354
rect 8962 -7698 9042 -7526
rect 8962 -7870 9042 -7698
rect 1170 -8278 1250 -8106
rect 3304 -8430 4006 -8368
rect 3304 -9010 3366 -8430
rect 3450 -8578 3858 -8518
rect 3450 -8868 3508 -8578
rect 3796 -8868 3858 -8578
rect 3450 -8922 3858 -8868
rect 3944 -9010 4006 -8430
rect 3304 -9072 4006 -9010
rect 4120 -8430 4822 -8368
rect 4120 -9010 4182 -8430
rect 4266 -8578 4674 -8518
rect 4266 -8868 4324 -8578
rect 4612 -8868 4674 -8578
rect 4266 -8922 4674 -8868
rect 4760 -9010 4822 -8430
rect 4120 -9072 4822 -9010
rect 4936 -8430 5638 -8368
rect 4936 -9010 4998 -8430
rect 5082 -8578 5490 -8518
rect 5082 -8868 5140 -8578
rect 5428 -8868 5490 -8578
rect 5082 -8922 5490 -8868
rect 5576 -9010 5638 -8430
rect 4936 -9072 5638 -9010
rect 5752 -8430 6454 -8368
rect 5752 -9010 5814 -8430
rect 5898 -8578 6306 -8518
rect 5898 -8868 5956 -8578
rect 6244 -8868 6306 -8578
rect 5898 -8922 6306 -8868
rect 6392 -9010 6454 -8430
rect 5752 -9072 6454 -9010
rect 6568 -8430 7270 -8368
rect 6568 -9010 6630 -8430
rect 6714 -8578 7122 -8518
rect 6714 -8868 6772 -8578
rect 7060 -8868 7122 -8578
rect 6714 -8922 7122 -8868
rect 7208 -9010 7270 -8430
rect 6568 -9072 7270 -9010
rect 3304 -9246 4006 -9184
rect 3304 -9826 3366 -9246
rect 3450 -9394 3858 -9334
rect 3450 -9684 3508 -9394
rect 3796 -9684 3858 -9394
rect 3450 -9738 3858 -9684
rect 3944 -9826 4006 -9246
rect 3304 -9888 4006 -9826
rect 4120 -9246 4822 -9184
rect 4120 -9826 4182 -9246
rect 4266 -9394 4674 -9334
rect 4266 -9684 4324 -9394
rect 4612 -9684 4674 -9394
rect 4266 -9738 4674 -9684
rect 4760 -9826 4822 -9246
rect 4120 -9888 4822 -9826
rect 4936 -9246 5638 -9184
rect 4936 -9826 4998 -9246
rect 5082 -9394 5490 -9334
rect 5082 -9684 5140 -9394
rect 5428 -9684 5490 -9394
rect 5082 -9738 5490 -9684
rect 5576 -9826 5638 -9246
rect 4936 -9888 5638 -9826
rect 5752 -9246 6454 -9184
rect 5752 -9826 5814 -9246
rect 5898 -9394 6306 -9334
rect 5898 -9684 5956 -9394
rect 6244 -9684 6306 -9394
rect 5898 -9738 6306 -9684
rect 6392 -9826 6454 -9246
rect 5752 -9888 6454 -9826
rect 6568 -9246 7270 -9184
rect 6568 -9826 6630 -9246
rect 6714 -9394 7122 -9334
rect 6714 -9684 6772 -9394
rect 7060 -9684 7122 -9394
rect 6714 -9738 7122 -9684
rect 7208 -9826 7270 -9246
rect 6568 -9888 7270 -9826
<< metal1 >>
rect 1960 -2488 2110 -2478
rect 1960 -2678 1972 -2488
rect 2100 -2678 2110 -2488
rect 1960 -2688 2110 -2678
rect 2390 -2488 2540 -2478
rect 2390 -2678 2402 -2488
rect 2530 -2678 2540 -2488
rect 1612 -3944 1684 -2800
rect 1988 -2812 2082 -2688
rect 1902 -3150 1954 -3144
rect 1902 -3412 1954 -3406
rect 1988 -3788 1994 -2812
rect 2028 -3788 2082 -2812
rect 2390 -2812 2540 -2678
rect 3454 -2488 3604 -2478
rect 3454 -2678 3466 -2488
rect 3594 -2678 3604 -2488
rect 2116 -3150 2168 -3144
rect 2116 -3412 2168 -3406
rect 1612 -4056 1620 -3944
rect 1676 -4056 1684 -3944
rect 1612 -5386 1684 -4056
rect 1724 -3838 1892 -3832
rect 1724 -4296 1892 -3890
rect 1724 -4354 1892 -4348
rect 1988 -4398 2082 -3788
rect 2390 -3788 2448 -2812
rect 2482 -3788 2540 -2812
rect 2172 -3838 2346 -3832
rect 2172 -3890 2178 -3838
rect 2172 -4296 2346 -3890
rect 2172 -4348 2178 -4296
rect 2172 -4354 2346 -4348
rect 1902 -4742 1954 -4736
rect 1902 -5004 1954 -4998
rect 1988 -5374 1994 -4398
rect 2028 -5374 2082 -4398
rect 2390 -4398 2540 -3788
rect 2942 -3832 3054 -2800
rect 3454 -2812 3604 -2678
rect 4518 -2488 4668 -2478
rect 4518 -2678 4530 -2488
rect 4658 -2678 4668 -2488
rect 3454 -3788 3512 -2812
rect 3546 -3788 3604 -2812
rect 2578 -3838 3416 -3832
rect 2578 -3890 2584 -3838
rect 2952 -3888 3042 -3838
rect 2952 -3890 2958 -3888
rect 2578 -3896 2958 -3890
rect 3036 -3890 3042 -3888
rect 3410 -3890 3416 -3838
rect 3036 -3896 3416 -3890
rect 2584 -4290 2952 -3896
rect 3042 -4290 3410 -3896
rect 2578 -4296 2958 -4290
rect 2578 -4348 2584 -4296
rect 2952 -4348 2958 -4296
rect 2578 -4354 2958 -4348
rect 3036 -4296 3416 -4290
rect 3036 -4348 3042 -4296
rect 3410 -4348 3416 -4296
rect 3036 -4354 3416 -4348
rect 2116 -4742 2168 -4736
rect 2116 -5004 2168 -4998
rect 1988 -5386 2082 -5374
rect 2390 -5374 2448 -4398
rect 2482 -5374 2540 -4398
rect 3454 -4398 3604 -3788
rect 4006 -3832 4118 -2800
rect 4518 -2812 4668 -2678
rect 4518 -3788 4576 -2812
rect 4610 -3788 4668 -2812
rect 5582 -2488 5732 -2478
rect 5582 -2678 5594 -2488
rect 5722 -2678 5732 -2488
rect 5582 -2812 5732 -2678
rect 5096 -2866 5154 -2860
rect 5096 -3784 5154 -3778
rect 3642 -3838 4480 -3832
rect 3642 -3890 3648 -3838
rect 4016 -3888 4106 -3838
rect 4016 -3890 4022 -3888
rect 3642 -3896 4022 -3890
rect 4100 -3890 4106 -3888
rect 4474 -3890 4480 -3838
rect 4100 -3896 4480 -3890
rect 3648 -4290 4016 -3896
rect 4106 -4290 4474 -3896
rect 3642 -4296 4022 -4290
rect 3642 -4348 3648 -4296
rect 4016 -4348 4022 -4296
rect 3642 -4354 4022 -4348
rect 4100 -4296 4480 -4290
rect 4100 -4348 4106 -4296
rect 4474 -4348 4480 -4296
rect 4100 -4354 4480 -4348
rect 2390 -5386 2540 -5374
rect 2968 -4464 3026 -4458
rect 2968 -5382 3026 -5376
rect 3454 -5374 3512 -4398
rect 3546 -5374 3604 -4398
rect 4518 -4398 4668 -3788
rect 5582 -3788 5640 -2812
rect 5674 -3788 5732 -2812
rect 6646 -2488 6796 -2478
rect 6646 -2678 6658 -2488
rect 6786 -2678 6796 -2488
rect 6646 -2812 6796 -2678
rect 4706 -3838 5086 -3832
rect 4706 -3890 4712 -3838
rect 5080 -3890 5086 -3838
rect 4706 -3896 5086 -3890
rect 5164 -3838 5544 -3832
rect 5164 -3890 5170 -3838
rect 5538 -3890 5544 -3838
rect 5164 -3896 5544 -3890
rect 4712 -4290 5080 -3896
rect 5170 -4290 5538 -3896
rect 4706 -4296 5544 -4290
rect 4706 -4348 4712 -4296
rect 5080 -4348 5170 -4296
rect 5538 -4348 5544 -4296
rect 4706 -4354 5544 -4348
rect 3454 -5386 3604 -5374
rect 4032 -4464 4090 -4458
rect 4032 -5382 4090 -5376
rect 4518 -5374 4576 -4398
rect 4610 -5374 4668 -4398
rect 4518 -5386 4668 -5374
rect 4958 -5830 5294 -4354
rect 5582 -4398 5732 -3788
rect 6160 -3412 6218 -3406
rect 6160 -3794 6218 -3788
rect 6646 -3788 6704 -2812
rect 6738 -3788 6796 -2812
rect 7892 -2486 7968 -2478
rect 7892 -2676 7898 -2486
rect 7962 -2676 7968 -2486
rect 5770 -3838 6150 -3832
rect 5770 -3890 5776 -3838
rect 6144 -3890 6150 -3838
rect 5770 -3896 6150 -3890
rect 6228 -3838 6608 -3832
rect 6228 -3890 6234 -3838
rect 6602 -3890 6608 -3838
rect 6228 -3896 6608 -3890
rect 5776 -4290 6144 -3896
rect 6234 -4290 6602 -3896
rect 5770 -4296 6150 -4290
rect 5770 -4348 5776 -4296
rect 6144 -4348 6150 -4296
rect 5770 -4354 6150 -4348
rect 6228 -4296 6608 -4290
rect 6228 -4348 6234 -4296
rect 6602 -4348 6608 -4296
rect 6228 -4354 6608 -4348
rect 5582 -5374 5640 -4398
rect 5674 -5374 5732 -4398
rect 6160 -4398 6218 -4392
rect 6160 -4780 6218 -4774
rect 6646 -4398 6796 -3788
rect 7224 -3412 7282 -3406
rect 7224 -3794 7282 -3788
rect 7354 -3410 7412 -3404
rect 7892 -3410 7968 -2676
rect 7354 -3792 7412 -3786
rect 7806 -3598 7864 -3588
rect 7806 -3794 7864 -3788
rect 7892 -3786 7898 -3410
rect 7932 -3786 7968 -3410
rect 7892 -3798 7968 -3786
rect 6834 -3838 7214 -3832
rect 6834 -3890 6840 -3838
rect 7208 -3890 7214 -3838
rect 6834 -3896 7214 -3890
rect 6840 -4290 7208 -3896
rect 7416 -3944 7808 -3884
rect 7416 -4056 7532 -3944
rect 7700 -4056 7808 -3944
rect 7416 -4068 7808 -4056
rect 7416 -4180 7532 -4068
rect 7700 -4180 7808 -4068
rect 6834 -4296 7214 -4290
rect 6834 -4348 6840 -4296
rect 7208 -4348 7214 -4296
rect 7416 -4300 7808 -4180
rect 6834 -4354 7214 -4348
rect 7912 -4386 7968 -3798
rect 8046 -3222 9480 -3156
rect 8046 -3944 8134 -3222
rect 9578 -3260 9634 -3248
rect 9492 -3568 9550 -3562
rect 9492 -3810 9550 -3804
rect 8046 -4180 8052 -3944
rect 8126 -4180 8134 -3944
rect 8046 -4186 8134 -4180
rect 9578 -4236 9584 -3260
rect 9618 -4236 9634 -3260
rect 8048 -4316 9480 -4312
rect 5582 -5386 5732 -5374
rect 6646 -5374 6704 -4398
rect 6738 -5374 6796 -4398
rect 7224 -4398 7282 -4392
rect 7224 -4780 7282 -4774
rect 7354 -4398 7412 -4392
rect 7806 -4398 7864 -4388
rect 7806 -4594 7864 -4588
rect 7892 -4398 7968 -4386
rect 7354 -4780 7412 -4774
rect 7892 -4774 7898 -4398
rect 7932 -4774 7968 -4398
rect 7892 -4786 7968 -4774
rect 8046 -4378 9480 -4316
rect 8046 -4724 8134 -4378
rect 9578 -4416 9634 -4236
rect 9578 -4442 9584 -4416
rect 8104 -4960 8134 -4724
rect 8046 -5342 8134 -4960
rect 6646 -5386 6796 -5374
rect 9504 -5392 9584 -4442
rect 9618 -4826 9634 -4416
rect 9618 -5392 9912 -4826
rect 9504 -5430 9912 -5392
rect 4958 -5962 4974 -5830
rect 5278 -5962 5294 -5830
rect 9166 -5476 9304 -5470
rect 9166 -5688 9172 -5476
rect 9298 -5688 9304 -5476
rect 4958 -6018 5294 -5962
rect 8956 -5978 9048 -5886
rect 1772 -6120 1778 -6064
rect 2146 -6120 2152 -6064
rect 2230 -6120 2236 -6064
rect 2604 -6120 2610 -6064
rect 2836 -6120 2842 -6064
rect 3210 -6120 3216 -6064
rect 3294 -6120 3300 -6064
rect 3668 -6120 3674 -6064
rect 3900 -6120 3906 -6064
rect 4274 -6120 4280 -6064
rect 4358 -6120 4364 -6064
rect 4732 -6120 4738 -6064
rect 5518 -6120 5524 -6064
rect 5892 -6120 5898 -6064
rect 6124 -6120 6130 -6064
rect 6498 -6120 6504 -6064
rect 6582 -6120 6588 -6064
rect 6956 -6120 6962 -6064
rect 7188 -6120 7194 -6064
rect 7562 -6120 7568 -6064
rect 7646 -6120 7652 -6064
rect 8020 -6120 8026 -6064
rect 8252 -6120 8258 -6064
rect 8626 -6120 8632 -6064
rect 1376 -7192 1514 -7186
rect 1146 -7418 1256 -7260
rect 1146 -8278 1170 -7418
rect 1250 -8278 1256 -7418
rect 1376 -7316 1382 -7192
rect 1508 -7316 1514 -7192
rect 1376 -7712 1514 -7316
rect 1636 -7350 1682 -6146
rect 1710 -7198 1766 -6192
rect 2162 -6206 2220 -6196
rect 2162 -7098 2220 -7088
rect 1710 -7316 1766 -7310
rect 2616 -7198 2672 -6192
rect 2616 -7316 2672 -7310
rect 2700 -7350 2746 -6146
rect 2774 -7198 2830 -6192
rect 3226 -6216 3284 -6206
rect 3226 -7108 3284 -7098
rect 2774 -7316 2830 -7310
rect 3680 -7198 3736 -6192
rect 3680 -7316 3736 -7310
rect 3764 -7350 3810 -6146
rect 3838 -7198 3894 -6192
rect 4290 -6216 4348 -6206
rect 4290 -7108 4348 -7098
rect 3838 -7316 3894 -7310
rect 4744 -7198 4800 -6192
rect 4744 -7316 4800 -7310
rect 4828 -7350 4874 -6146
rect 5988 -6158 6034 -6146
rect 5450 -6218 5508 -6208
rect 5450 -7110 5508 -7100
rect 5220 -7184 5354 -7176
rect 5220 -7308 5228 -7184
rect 5348 -7308 5354 -7184
rect 5904 -7190 5960 -6198
rect 5904 -7308 5960 -7302
rect 5988 -7134 5994 -6158
rect 6028 -7134 6034 -6158
rect 7052 -6158 7098 -6146
rect 1632 -7356 1804 -7350
rect 1686 -7456 1804 -7356
rect 1146 -10132 1256 -8278
rect 1146 -10564 1170 -10132
rect 1250 -10564 1256 -10132
rect 1146 -10574 1256 -10564
rect 1632 -10136 1804 -7456
rect 2696 -7356 2750 -7350
rect 2696 -7462 2750 -7456
rect 3760 -7356 3814 -7350
rect 3760 -7462 3814 -7456
rect 4824 -7356 4878 -7350
rect 4824 -7462 4878 -7456
rect 5220 -7680 5354 -7308
rect 5988 -7350 6034 -7134
rect 6062 -7190 6118 -6198
rect 6514 -6218 6572 -6208
rect 6514 -7110 6572 -7100
rect 6062 -7308 6118 -7302
rect 6968 -7190 7024 -6198
rect 6968 -7308 7024 -7302
rect 7052 -7134 7058 -6158
rect 7092 -7134 7098 -6158
rect 8116 -6158 8162 -6146
rect 7052 -7350 7098 -7134
rect 7126 -7190 7182 -6198
rect 7578 -6218 7636 -6208
rect 7578 -7110 7636 -7100
rect 7126 -7308 7182 -7302
rect 8032 -7190 8088 -6198
rect 8032 -7308 8088 -7302
rect 8116 -7134 8122 -6158
rect 8156 -7134 8162 -6158
rect 8116 -7350 8162 -7134
rect 8190 -7190 8246 -6198
rect 8642 -6218 8700 -6208
rect 8642 -7110 8700 -7100
rect 8956 -7146 8962 -5978
rect 8190 -7308 8246 -7302
rect 5984 -7356 6038 -7350
rect 5984 -7462 6038 -7456
rect 7048 -7356 7102 -7350
rect 7048 -7462 7102 -7456
rect 8112 -7356 8166 -7350
rect 8112 -7462 8166 -7456
rect 5218 -7690 5358 -7680
rect 5218 -7814 5228 -7690
rect 5348 -7814 5358 -7690
rect 5218 -7822 5358 -7814
rect 8938 -7870 8962 -7146
rect 9042 -7870 9048 -5978
rect 9166 -6122 9304 -5688
rect 9792 -7360 9912 -5430
rect 9986 -5476 10238 -4936
rect 9986 -5688 10048 -5476
rect 10174 -5688 10238 -5476
rect 9986 -6230 10238 -5688
rect 9792 -7452 9800 -7360
rect 9904 -7452 9912 -7360
rect 1632 -10568 1638 -10136
rect 1798 -10568 1804 -10136
rect 1632 -10574 1804 -10568
rect 3294 -8368 7276 -8354
rect 3294 -9072 3304 -8368
rect 3366 -8518 3944 -8430
rect 3366 -8922 3450 -8518
rect 3508 -8584 3796 -8578
rect 3508 -8862 3514 -8584
rect 3588 -8654 3720 -8646
rect 3588 -8794 3720 -8786
rect 3790 -8862 3796 -8584
rect 3508 -8868 3796 -8862
rect 3858 -8922 3944 -8518
rect 3366 -9010 3944 -8922
rect 4006 -8886 4120 -8368
rect 4006 -9072 4012 -8886
rect 3294 -9088 4012 -9072
rect 4110 -9072 4120 -8886
rect 4182 -8518 4760 -8430
rect 4182 -8922 4266 -8518
rect 4324 -8584 4612 -8578
rect 4324 -8862 4330 -8584
rect 4404 -8654 4536 -8646
rect 4404 -8794 4536 -8786
rect 4606 -8862 4612 -8584
rect 4324 -8868 4612 -8862
rect 4674 -8922 4760 -8518
rect 4182 -9010 4760 -8922
rect 4822 -8886 4936 -8368
rect 4822 -9072 4828 -8886
rect 4110 -9088 4828 -9072
rect 4926 -9072 4936 -8886
rect 4998 -8518 5576 -8430
rect 4998 -8922 5082 -8518
rect 5140 -8584 5428 -8578
rect 5140 -8862 5146 -8584
rect 5220 -8654 5352 -8646
rect 5220 -8794 5352 -8786
rect 5422 -8862 5428 -8584
rect 5140 -8868 5428 -8862
rect 5490 -8922 5576 -8518
rect 4998 -9010 5576 -8922
rect 5638 -8886 5752 -8368
rect 5638 -9072 5644 -8886
rect 4926 -9088 5644 -9072
rect 5742 -9072 5752 -8886
rect 5814 -8518 6392 -8430
rect 5814 -8922 5898 -8518
rect 5956 -8584 6244 -8578
rect 5956 -8862 5962 -8584
rect 6036 -8654 6168 -8646
rect 6036 -8794 6168 -8786
rect 6238 -8862 6244 -8584
rect 5956 -8868 6244 -8862
rect 6306 -8922 6392 -8518
rect 5814 -9010 6392 -8922
rect 6454 -8884 6568 -8368
rect 6454 -9072 6460 -8884
rect 5742 -9088 6460 -9072
rect 6558 -9072 6568 -8884
rect 6630 -8518 7208 -8430
rect 6630 -8922 6714 -8518
rect 6772 -8584 7060 -8578
rect 6772 -8862 6778 -8584
rect 6852 -8654 6984 -8646
rect 6852 -8794 6984 -8786
rect 7054 -8862 7060 -8584
rect 6772 -8868 7060 -8862
rect 7122 -8922 7208 -8518
rect 6630 -9010 7208 -8922
rect 7270 -9072 7276 -8368
rect 6558 -9088 7276 -9072
rect 3294 -9170 3822 -9088
rect 6758 -9170 7276 -9088
rect 3294 -9184 4012 -9170
rect 3294 -9888 3304 -9184
rect 3366 -9334 3944 -9246
rect 3366 -9738 3450 -9334
rect 3508 -9402 3796 -9394
rect 3508 -9678 3514 -9402
rect 3588 -9470 3720 -9462
rect 3588 -9610 3720 -9602
rect 3790 -9678 3796 -9402
rect 3508 -9684 3796 -9678
rect 3858 -9738 3944 -9334
rect 3366 -9826 3944 -9738
rect 4006 -9366 4012 -9184
rect 4110 -9184 4828 -9170
rect 4110 -9366 4120 -9184
rect 4006 -9888 4120 -9366
rect 4182 -9334 4760 -9246
rect 4182 -9738 4266 -9334
rect 4324 -9400 4612 -9394
rect 4324 -9678 4330 -9400
rect 4404 -9470 4536 -9462
rect 4404 -9610 4536 -9602
rect 4606 -9678 4612 -9400
rect 4324 -9684 4612 -9678
rect 4674 -9738 4760 -9334
rect 4182 -9826 4760 -9738
rect 4822 -9366 4828 -9184
rect 4926 -9184 5644 -9170
rect 4926 -9366 4936 -9184
rect 4822 -9888 4936 -9366
rect 4998 -9334 5576 -9246
rect 4998 -9738 5082 -9334
rect 5140 -9400 5428 -9394
rect 5140 -9678 5146 -9400
rect 5220 -9470 5352 -9462
rect 5220 -9610 5352 -9602
rect 5422 -9678 5428 -9400
rect 5140 -9684 5428 -9678
rect 5490 -9738 5576 -9334
rect 4998 -9826 5576 -9738
rect 5638 -9366 5644 -9184
rect 5742 -9184 6460 -9170
rect 5742 -9366 5752 -9184
rect 5638 -9888 5752 -9366
rect 5814 -9334 6392 -9246
rect 5814 -9738 5898 -9334
rect 5956 -9400 6244 -9394
rect 5956 -9678 5962 -9400
rect 6036 -9470 6168 -9462
rect 6036 -9610 6168 -9602
rect 6238 -9678 6244 -9400
rect 5956 -9684 6244 -9678
rect 6306 -9738 6392 -9334
rect 5814 -9826 6392 -9738
rect 6454 -9366 6460 -9184
rect 6558 -9184 7276 -9170
rect 6558 -9366 6568 -9184
rect 6454 -9888 6568 -9366
rect 6630 -9334 7208 -9246
rect 6630 -9738 6714 -9334
rect 6772 -9400 7060 -9394
rect 6772 -9678 6778 -9400
rect 6852 -9470 6984 -9462
rect 6852 -9610 6984 -9602
rect 7054 -9678 7060 -9400
rect 6772 -9684 7060 -9678
rect 7122 -9738 7208 -9334
rect 6630 -9826 7208 -9738
rect 7270 -9888 7276 -9184
rect 3294 -9904 7276 -9888
rect 3294 -10148 4868 -9904
rect 3294 -10540 3314 -10148
rect 4842 -10540 4868 -10148
rect 3294 -10574 4868 -10540
rect 5700 -10150 7274 -9904
rect 5700 -10542 5720 -10150
rect 7248 -10542 7274 -10150
rect 5700 -10574 7274 -10542
rect 8938 -10132 9048 -7870
rect 9166 -9966 9304 -7864
rect 9166 -10076 9178 -9966
rect 9294 -10076 9304 -9966
rect 9166 -10088 9304 -10076
rect 8938 -10564 8952 -10132
rect 9032 -10564 9048 -10132
rect 8938 -10574 9048 -10564
rect 9792 -10132 9912 -7452
rect 9792 -10564 9810 -10132
rect 9890 -10564 9912 -10132
rect 9792 -10574 9912 -10564
<< via1 >>
rect 1972 -2678 2100 -2488
rect 2402 -2678 2530 -2488
rect 1902 -3406 1954 -3150
rect 3466 -2678 3594 -2488
rect 2116 -3406 2168 -3150
rect 1620 -4056 1676 -3944
rect 1724 -3890 1892 -3838
rect 1724 -4348 1892 -4296
rect 2178 -3890 2346 -3838
rect 2178 -4348 2346 -4296
rect 1902 -4998 1954 -4742
rect 4530 -2678 4658 -2488
rect 2584 -3890 2952 -3838
rect 3042 -3890 3410 -3838
rect 2584 -4348 2952 -4296
rect 3042 -4348 3410 -4296
rect 2116 -4998 2168 -4742
rect 5594 -2678 5722 -2488
rect 5096 -3778 5154 -2866
rect 3648 -3890 4016 -3838
rect 4106 -3890 4474 -3838
rect 3648 -4348 4016 -4296
rect 4106 -4348 4474 -4296
rect 2968 -5376 3026 -4464
rect 6658 -2678 6786 -2488
rect 4712 -3890 5080 -3838
rect 5170 -3890 5538 -3838
rect 4712 -4348 5080 -4296
rect 5170 -4348 5538 -4296
rect 4032 -5376 4090 -4464
rect 6160 -3788 6218 -3412
rect 7898 -2676 7962 -2486
rect 5776 -3890 6144 -3838
rect 6234 -3890 6602 -3838
rect 5776 -4348 6144 -4296
rect 6234 -4348 6602 -4296
rect 6160 -4774 6218 -4398
rect 7224 -3788 7282 -3412
rect 7354 -3786 7412 -3410
rect 7806 -3788 7864 -3598
rect 6840 -3890 7208 -3838
rect 7532 -4056 7700 -3944
rect 7532 -4180 7700 -4068
rect 6840 -4348 7208 -4296
rect 9492 -3804 9550 -3568
rect 8052 -4180 8126 -3944
rect 7224 -4774 7282 -4398
rect 7354 -4774 7412 -4398
rect 7806 -4588 7864 -4398
rect 8046 -4960 8104 -4724
rect 4974 -5962 5278 -5830
rect 9172 -5688 9298 -5476
rect 1778 -6120 2146 -6064
rect 2236 -6120 2604 -6064
rect 2842 -6120 3210 -6064
rect 3300 -6120 3668 -6064
rect 3906 -6120 4274 -6064
rect 4364 -6120 4732 -6064
rect 5524 -6120 5892 -6064
rect 6130 -6120 6498 -6064
rect 6588 -6120 6956 -6064
rect 7194 -6120 7562 -6064
rect 7652 -6120 8020 -6064
rect 8258 -6120 8626 -6064
rect 1382 -7316 1508 -7192
rect 2162 -7088 2220 -6206
rect 1710 -7310 1766 -7198
rect 2616 -7310 2672 -7198
rect 3226 -7098 3284 -6216
rect 2774 -7310 2830 -7198
rect 3680 -7310 3736 -7198
rect 4290 -7098 4348 -6216
rect 3838 -7310 3894 -7198
rect 4744 -7310 4800 -7198
rect 5450 -7100 5508 -6218
rect 5228 -7308 5348 -7184
rect 5904 -7302 5960 -7190
rect 1632 -7456 1686 -7356
rect 1392 -8192 1498 -7968
rect 1170 -10564 1250 -10132
rect 2696 -7456 2750 -7356
rect 3760 -7456 3814 -7356
rect 4824 -7456 4878 -7356
rect 6514 -7100 6572 -6218
rect 6062 -7302 6118 -7190
rect 6968 -7302 7024 -7190
rect 7578 -7100 7636 -6218
rect 7126 -7302 7182 -7190
rect 8032 -7302 8088 -7190
rect 8642 -7100 8700 -6218
rect 8190 -7302 8246 -7190
rect 5984 -7456 6038 -7356
rect 7048 -7456 7102 -7356
rect 8112 -7456 8166 -7356
rect 5228 -7814 5348 -7690
rect 10048 -5688 10174 -5476
rect 9800 -7452 9904 -7360
rect 1638 -10568 1798 -10136
rect 3588 -8786 3720 -8654
rect 4404 -8786 4536 -8654
rect 5220 -8786 5352 -8654
rect 6036 -8786 6168 -8654
rect 6852 -8786 6984 -8654
rect 3588 -9602 3720 -9470
rect 4404 -9602 4536 -9470
rect 5220 -9602 5352 -9470
rect 6036 -9602 6168 -9470
rect 6852 -9602 6984 -9470
rect 3314 -10540 4842 -10148
rect 5720 -10542 7248 -10150
rect 9178 -10076 9294 -9966
rect 8952 -10564 9032 -10132
rect 9810 -10564 9890 -10132
<< metal2 >>
rect 1044 -2486 10268 -2240
rect 1044 -2488 7898 -2486
rect 1044 -2678 1972 -2488
rect 2100 -2678 2402 -2488
rect 2530 -2678 3466 -2488
rect 3594 -2678 4530 -2488
rect 4658 -2678 5594 -2488
rect 5722 -2678 6658 -2488
rect 6786 -2676 7898 -2488
rect 7962 -2676 10268 -2486
rect 6786 -2678 10268 -2676
rect 1044 -2688 10268 -2678
rect 5096 -2866 5154 -2856
rect 1902 -3150 2168 -3140
rect 1964 -3406 2106 -3150
rect 1902 -3416 2168 -3406
rect 5096 -3788 5154 -3778
rect 6160 -3410 7412 -3400
rect 6160 -3412 7354 -3410
rect 6218 -3788 7224 -3412
rect 7282 -3786 7354 -3412
rect 8718 -3568 9550 -3562
rect 7282 -3788 7412 -3786
rect 6160 -3798 7412 -3788
rect 7806 -3598 7864 -3588
rect 7806 -3798 7864 -3788
rect 8718 -3804 9492 -3568
rect 8718 -3810 9550 -3804
rect 1718 -3834 7874 -3826
rect 1718 -3838 7806 -3834
rect 1718 -3890 1724 -3838
rect 1892 -3890 2178 -3838
rect 2346 -3890 2584 -3838
rect 2952 -3890 3042 -3838
rect 3410 -3890 3648 -3838
rect 4016 -3890 4106 -3838
rect 4474 -3890 4712 -3838
rect 5080 -3890 5170 -3838
rect 5538 -3890 5776 -3838
rect 6144 -3890 6234 -3838
rect 6602 -3890 6840 -3838
rect 7208 -3890 7806 -3838
rect 7864 -3890 7874 -3834
rect 1718 -3902 7874 -3890
rect 1614 -3944 8132 -3938
rect 1614 -4056 1620 -3944
rect 1676 -4056 7532 -3944
rect 7700 -4056 8052 -3944
rect 1614 -4062 8052 -4056
rect 7532 -4068 8052 -4062
rect 7700 -4180 8052 -4068
rect 8126 -4180 8132 -3944
rect 7532 -4186 8132 -4180
rect 1718 -4292 7874 -4284
rect 1718 -4296 7806 -4292
rect 1718 -4348 1724 -4296
rect 1892 -4348 2178 -4296
rect 2346 -4348 2584 -4296
rect 2952 -4348 3042 -4296
rect 3410 -4348 3648 -4296
rect 4016 -4348 4106 -4296
rect 4474 -4348 4712 -4296
rect 5080 -4348 5170 -4296
rect 5538 -4348 5776 -4296
rect 6144 -4348 6234 -4296
rect 6602 -4348 6840 -4296
rect 7208 -4348 7806 -4296
rect 7864 -4348 7874 -4292
rect 1718 -4360 7874 -4348
rect 6160 -4398 7412 -4388
rect 2968 -4464 3026 -4454
rect 1902 -4742 2168 -4732
rect 1964 -4998 2106 -4742
rect 1902 -5008 2168 -4998
rect 2936 -5376 2968 -5324
rect 4032 -4464 4090 -4454
rect 3026 -5376 3056 -5324
rect 2936 -5470 3056 -5376
rect 4000 -5376 4032 -5324
rect 6218 -4774 7224 -4398
rect 7282 -4774 7354 -4398
rect 7806 -4398 7864 -4388
rect 7806 -4598 7864 -4588
rect 8718 -4718 8966 -3810
rect 6160 -4786 7412 -4774
rect 8040 -4724 8966 -4718
rect 8040 -4960 8046 -4724
rect 8104 -4960 8966 -4724
rect 8040 -4966 8966 -4960
rect 4090 -5376 4120 -5324
rect 4000 -5470 4120 -5376
rect 2936 -5476 10238 -5470
rect 2936 -5688 9172 -5476
rect 9298 -5688 10048 -5476
rect 10174 -5688 10238 -5476
rect 2936 -5694 10238 -5688
rect 4974 -5830 5278 -5820
rect 4974 -5972 5278 -5962
rect 1772 -6064 8700 -6054
rect 1772 -6120 1778 -6064
rect 2146 -6120 2236 -6064
rect 2604 -6120 2842 -6064
rect 3210 -6120 3300 -6064
rect 3668 -6120 3906 -6064
rect 4274 -6120 4364 -6064
rect 4732 -6120 5524 -6064
rect 5892 -6120 6130 -6064
rect 6498 -6120 6588 -6064
rect 6956 -6120 7194 -6064
rect 7562 -6120 7652 -6064
rect 8020 -6120 8258 -6064
rect 8626 -6120 8700 -6064
rect 1772 -6130 8700 -6120
rect 2162 -6206 2220 -6196
rect 2162 -7098 2220 -7088
rect 3226 -6216 3284 -6206
rect 3226 -7108 3284 -7098
rect 4290 -6216 4348 -6206
rect 4290 -7108 4348 -7098
rect 5450 -6218 5508 -6130
rect 5450 -7110 5508 -7100
rect 6514 -6218 6572 -6130
rect 6514 -7110 6572 -7100
rect 7578 -6218 7636 -6130
rect 7578 -7110 7636 -7100
rect 8642 -6218 8700 -6130
rect 8642 -7110 8700 -7100
rect 5220 -7184 8246 -7176
rect 1376 -7192 4800 -7186
rect 1376 -7316 1382 -7192
rect 1508 -7198 4800 -7192
rect 1508 -7310 1710 -7198
rect 1766 -7310 2616 -7198
rect 2672 -7310 2774 -7198
rect 2830 -7310 3680 -7198
rect 3736 -7310 3838 -7198
rect 3894 -7310 4744 -7198
rect 1508 -7316 4800 -7310
rect 5220 -7308 5228 -7184
rect 5348 -7190 8246 -7184
rect 5348 -7302 5904 -7190
rect 5960 -7302 6062 -7190
rect 6118 -7302 6968 -7190
rect 7024 -7302 7126 -7190
rect 7182 -7302 8032 -7190
rect 8088 -7302 8190 -7190
rect 5348 -7308 8246 -7302
rect 5220 -7316 8246 -7308
rect 1376 -7322 4800 -7316
rect 1632 -7356 9912 -7350
rect 1686 -7456 2696 -7356
rect 2750 -7456 3760 -7356
rect 3814 -7456 4824 -7356
rect 4878 -7456 5984 -7356
rect 6038 -7456 7048 -7356
rect 7102 -7456 8112 -7356
rect 8166 -7360 9912 -7356
rect 8166 -7452 9800 -7360
rect 9904 -7452 9912 -7360
rect 8166 -7456 9912 -7452
rect 1632 -7462 9912 -7456
rect 5218 -7690 5358 -7680
rect 5218 -7814 5228 -7690
rect 5348 -7814 5358 -7690
rect 5218 -7822 5358 -7814
rect 1392 -7968 6984 -7962
rect 1498 -8192 6984 -7968
rect 1392 -8198 6984 -8192
rect 3588 -8646 3720 -8198
rect 4404 -8646 4536 -8198
rect 3588 -8654 4536 -8646
rect 3720 -8786 4404 -8654
rect 3588 -8794 4536 -8786
rect 5220 -8654 5352 -8646
rect 5220 -8794 5352 -8786
rect 6036 -8654 6168 -8198
rect 6852 -8654 6984 -8198
rect 6168 -8786 6852 -8654
rect 6036 -8794 6984 -8786
rect 3588 -9462 3720 -8794
rect 4404 -9462 4536 -8794
rect 3588 -9470 4536 -9462
rect 3720 -9602 4404 -9470
rect 3588 -9610 4536 -9602
rect 5220 -9470 5352 -9462
rect 5220 -9956 5352 -9602
rect 6036 -9470 6168 -8794
rect 6852 -9470 6984 -8794
rect 6168 -9602 6852 -9470
rect 6036 -9610 6984 -9602
rect 5220 -9966 9304 -9956
rect 5220 -10076 9178 -9966
rect 9294 -10076 9304 -9966
rect 5220 -10088 9304 -10076
rect 1044 -10132 10268 -10126
rect 1044 -10564 1170 -10132
rect 1250 -10136 8952 -10132
rect 1250 -10564 1638 -10136
rect 1044 -10568 1638 -10564
rect 1798 -10148 8952 -10136
rect 1798 -10540 3314 -10148
rect 4842 -10150 8952 -10148
rect 4842 -10540 5720 -10150
rect 1798 -10542 5720 -10540
rect 7248 -10542 8952 -10150
rect 1798 -10564 8952 -10542
rect 9032 -10564 9810 -10132
rect 9890 -10564 10268 -10132
rect 1798 -10568 10268 -10564
rect 1044 -10574 10268 -10568
<< via2 >>
rect 1908 -3406 1954 -3150
rect 1954 -3406 1964 -3150
rect 2106 -3406 2116 -3150
rect 2116 -3406 2162 -3150
rect 5096 -3778 5154 -2866
rect 6160 -3788 6218 -3412
rect 7224 -3788 7282 -3412
rect 7354 -3786 7412 -3410
rect 7806 -3788 7864 -3598
rect 7806 -3890 7864 -3834
rect 7806 -4348 7864 -4292
rect 1908 -4998 1954 -4742
rect 1954 -4998 1964 -4742
rect 2106 -4998 2116 -4742
rect 2116 -4998 2162 -4742
rect 2968 -5376 3026 -4464
rect 4032 -5376 4090 -4464
rect 6160 -4774 6218 -4398
rect 7224 -4774 7282 -4398
rect 7354 -4774 7412 -4398
rect 7806 -4588 7864 -4398
rect 4974 -5962 5278 -5830
rect 2162 -7088 2220 -6206
rect 3226 -7098 3284 -6216
rect 4290 -7098 4348 -6216
rect 5450 -7100 5508 -6218
rect 6514 -7100 6572 -6218
rect 7578 -7100 7636 -6218
rect 8642 -7100 8700 -6218
rect 5228 -7814 5348 -7690
rect 5228 -8784 5344 -8662
<< metal3 >>
rect 5064 -2866 5184 -2856
rect 1902 -3150 2168 -3140
rect 1902 -3406 1908 -3150
rect 1964 -3406 2106 -3150
rect 2162 -3406 2168 -3150
rect 1902 -4742 2168 -3406
rect 5064 -3778 5096 -2866
rect 5154 -3778 5184 -2866
rect 1902 -4998 1908 -4742
rect 1964 -4998 2106 -4742
rect 2162 -4998 2168 -4742
rect 1902 -5008 2168 -4998
rect 2936 -4132 3056 -4128
rect 2936 -4244 2966 -4132
rect 3030 -4244 3056 -4132
rect 2936 -4464 3056 -4244
rect 2936 -5376 2968 -4464
rect 3026 -5376 3056 -4464
rect 2936 -5386 3056 -5376
rect 4000 -4132 4120 -4128
rect 4000 -4244 4030 -4132
rect 4094 -4244 4120 -4132
rect 4000 -4464 4120 -4244
rect 5064 -4132 5184 -3778
rect 5064 -4244 5094 -4132
rect 5158 -4244 5184 -4132
rect 5064 -4248 5184 -4244
rect 6128 -3412 6248 -3400
rect 6128 -3788 6160 -3412
rect 6218 -3788 6248 -3412
rect 4000 -5376 4032 -4464
rect 4090 -5376 4120 -4464
rect 4000 -5386 4120 -5376
rect 6128 -4398 6248 -3788
rect 6128 -4774 6160 -4398
rect 6218 -4774 6248 -4398
rect 6128 -5778 6248 -4774
rect 7218 -3410 7418 -3398
rect 7218 -3412 7354 -3410
rect 7218 -3788 7224 -3412
rect 7282 -3786 7354 -3412
rect 7412 -3786 7418 -3410
rect 7282 -3788 7418 -3786
rect 7218 -4398 7418 -3788
rect 7218 -4774 7224 -4398
rect 7282 -4774 7354 -4398
rect 7412 -4774 7418 -4398
rect 7796 -3598 7874 -3588
rect 7796 -3788 7806 -3598
rect 7864 -3788 7874 -3598
rect 7796 -3834 7874 -3788
rect 7796 -3890 7806 -3834
rect 7864 -3890 7874 -3834
rect 7796 -4292 7874 -3890
rect 7796 -4348 7806 -4292
rect 7864 -4348 7874 -4292
rect 7796 -4398 7874 -4348
rect 7796 -4588 7806 -4398
rect 7864 -4588 7874 -4398
rect 7796 -4598 7874 -4588
rect 7218 -5778 7418 -4774
rect 2132 -5830 5294 -5778
rect 2132 -5962 4974 -5830
rect 5278 -5962 5294 -5830
rect 2132 -6018 5294 -5962
rect 5420 -6018 8732 -5778
rect 2132 -6206 2252 -6018
rect 2132 -7088 2162 -6206
rect 2220 -7088 2252 -6206
rect 2132 -7098 2252 -7088
rect 3196 -6216 3316 -6018
rect 3196 -7098 3226 -6216
rect 3284 -7098 3316 -6216
rect 3196 -7108 3316 -7098
rect 4260 -6216 4380 -6018
rect 4260 -7098 4290 -6216
rect 4348 -7098 4380 -6216
rect 4260 -7108 4380 -7098
rect 5420 -6218 5540 -6018
rect 5420 -7100 5450 -6218
rect 5508 -7100 5540 -6218
rect 5420 -7110 5540 -7100
rect 6484 -6218 6604 -6018
rect 6484 -7100 6514 -6218
rect 6572 -7100 6604 -6218
rect 6484 -7110 6604 -7100
rect 7548 -6218 7668 -6018
rect 7548 -7100 7578 -6218
rect 7636 -7100 7668 -6218
rect 7548 -7110 7668 -7100
rect 8612 -6218 8732 -6018
rect 8612 -7100 8642 -6218
rect 8700 -7100 8732 -6218
rect 8612 -7110 8732 -7100
rect 5218 -7690 5358 -7680
rect 5218 -7814 5228 -7690
rect 5348 -7814 5358 -7690
rect 5218 -7822 5358 -7814
rect 5220 -8662 5352 -8646
rect 5220 -8784 5228 -8662
rect 5344 -8784 5352 -8662
rect 5220 -8794 5352 -8784
<< via3 >>
rect 2966 -4244 3030 -4132
rect 4030 -4244 4094 -4132
rect 5094 -4244 5158 -4132
rect 5228 -7814 5348 -7690
rect 5228 -8784 5344 -8662
<< metal4 >>
rect 2936 -4132 5184 -4128
rect 2936 -4244 2966 -4132
rect 3030 -4244 4030 -4132
rect 4094 -4244 5094 -4132
rect 5158 -4244 5184 -4132
rect 2936 -4248 5184 -4244
rect 5218 -7690 5358 -7680
rect 5218 -7814 5228 -7690
rect 5348 -7814 5358 -7690
rect 5218 -7822 5358 -7814
rect 5220 -8662 5352 -7822
rect 5220 -8784 5228 -8662
rect 5344 -8784 5352 -8662
rect 5220 -8794 5352 -8784
use sky130_fd_pr__nfet_01v8_lvt_69LV2L  M1
timestamp 1681576725
transform -1 0 8798 0 1 -3717
box -758 -557 758 557
use sky130_fd_pr__nfet_01v8_lvt_69LV2L  M2
timestamp 1681576725
transform -1 0 8798 0 1 -4873
box -758 -557 758 557
use sky130_fd_pr__pfet_01v8_lvt_SF68ZM  M31
timestamp 1681400668
transform -1 0 1808 0 1 -3336
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_SPM7ZP  M32
timestamp 1681402674
transform -1 0 1808 0 1 -4850
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_SF68ZM  M41
timestamp 1681400668
transform -1 0 2262 0 1 -3336
box -194 -564 194 598
use sky130_fd_pr__pfet_01v8_lvt_SPM7ZP  M42
timestamp 1681402674
transform -1 0 2262 0 1 -4850
box -194 -598 194 564
use sky130_fd_pr__pfet_01v8_lvt_HLVWZV  M51
timestamp 1681405906
transform -1 0 7612 0 1 -3634
box -294 -264 294 298
use sky130_fd_pr__pfet_01v8_lvt_MEMUZX  M52
timestamp 1681405906
transform -1 0 7612 0 1 -4550
box -294 -298 294 264
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M61
timestamp 1681402674
transform 1 0 5960 0 1 -3336
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M62
timestamp 1681402674
transform -1 0 6418 0 1 -3336
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M63
timestamp 1681402674
transform 1 0 7024 0 1 -3336
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M64
timestamp 1681402674
transform 1 0 5960 0 1 -4850
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M65
timestamp 1681402674
transform -1 0 6418 0 1 -4850
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M66
timestamp 1681402674
transform 1 0 7024 0 1 -4850
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M71
timestamp 1681402674
transform 1 0 2768 0 1 -3336
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M72
timestamp 1681402674
transform -1 0 3226 0 1 -3336
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M73
timestamp 1681402674
transform 1 0 3832 0 1 -3336
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M74
timestamp 1681402674
transform -1 0 4290 0 1 -3336
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M75
timestamp 1681402674
transform 1 0 4896 0 1 -4850
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M76
timestamp 1681402674
transform -1 0 5354 0 1 -4850
box -294 -598 294 564
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M81
timestamp 1681505393
transform -1 0 5708 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M82
timestamp 1681505393
transform 1 0 6314 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M83
timestamp 1681505393
transform -1 0 6772 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M84
timestamp 1681505393
transform 1 0 7378 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M85
timestamp 1681505393
transform -1 0 7836 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M86
timestamp 1681505393
transform 1 0 8442 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M91
timestamp 1681505393
transform 1 0 1962 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M92
timestamp 1681505393
transform -1 0 2420 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M93
timestamp 1681505393
transform 1 0 3026 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M94
timestamp 1681505393
transform -1 0 3484 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M95
timestamp 1681505393
transform 1 0 4090 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_D8YEEC  M96
timestamp 1681505393
transform -1 0 4548 0 1 -6615
box -258 -557 258 557
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M101
timestamp 1681402674
transform 1 0 4896 0 1 -3336
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M102
timestamp 1681402674
transform -1 0 5354 0 1 -3336
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M103
timestamp 1681402674
transform 1 0 2768 0 1 -4850
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M104
timestamp 1681402674
transform -1 0 3226 0 1 -4850
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M105
timestamp 1681402674
transform 1 0 3832 0 1 -4850
box -294 -598 294 564
use sky130_fd_pr__pfet_01v8_lvt_ME68ZX  M106
timestamp 1681402674
transform -1 0 4290 0 1 -4850
box -294 -598 294 564
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q1 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1671677353
transform 1 0 4888 0 1 -9118
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q3
timestamp 1671677353
transform 1 0 4888 0 1 -9934
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q21
timestamp 1671677353
transform 1 0 4072 0 1 -9118
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q22
timestamp 1671677353
transform 1 0 4072 0 1 -9934
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q23
timestamp 1671677353
transform 1 0 3256 0 1 -9118
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q24
timestamp 1671677353
transform 1 0 3256 0 1 -9934
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q25
timestamp 1671677353
transform 1 0 5704 0 1 -9118
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q26
timestamp 1671677353
transform 1 0 5704 0 1 -9934
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q27
timestamp 1671677353
transform 1 0 6520 0 1 -9118
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q28
timestamp 1671677353
transform 1 0 6520 0 1 -9934
box 0 0 796 796
use sky130_fd_pr__res_xhigh_po_0p69_7QK33H  XR3
timestamp 1680257378
transform 1 0 1445 0 1 -7786
box -71 -526 71 526
use sky130_fd_pr__res_xhigh_po_0p69_MTJZ47  XR4
timestamp 1680257378
transform 1 0 9235 0 1 -6918
box -71 -1032 71 1032
<< labels >>
flabel metal1 9986 -6230 10238 -4936 0 FreeMono 1600 90 0 0 out
port 2 nsew
flabel metal2 1044 -10574 10268 -10126 0 FreeMono 2400 0 0 0 vss
port 1 nsew
flabel metal2 1044 -2688 10268 -2240 0 FreeMono 2400 0 0 0 vdd
port 0 nsew
<< end >>
