magic
tech sky130A
timestamp 1682257739
<< metal1 >>
rect 136996 44211 145732 44214
rect 136996 43983 136999 44211
rect 137227 43983 145501 44211
rect 145729 43983 145732 44211
rect 136996 43980 145732 43983
rect 137444 38791 137844 38832
rect 138058 36275 138340 36313
rect 138058 36241 138390 36275
rect 138058 35681 138699 36241
rect 136164 35602 137230 35607
rect 136164 35379 136169 35602
rect 136392 35601 137230 35602
rect 136392 35379 137002 35601
rect 136164 35378 137002 35379
rect 137225 35378 137230 35601
rect 138058 35430 138102 35681
rect 138671 35430 138699 35681
rect 138058 35425 138699 35430
rect 136164 35373 137230 35378
rect 149309 23744 149703 23838
rect 137470 23739 149703 23744
rect 137470 23249 149355 23739
rect 149698 23249 149703 23739
rect 137470 23244 149703 23249
rect 149309 23155 149703 23244
rect 149309 23154 149684 23155
rect 137470 22923 139709 22928
rect 137470 22433 139309 22923
rect 139704 22433 139709 22923
rect 137470 22428 139709 22433
<< via1 >>
rect 136999 43983 137227 44211
rect 145501 43983 145729 44211
rect 136169 35379 136392 35602
rect 137002 35378 137225 35601
rect 138102 35430 138671 35681
rect 149355 23249 149698 23739
rect 139309 22433 139704 22923
<< metal2 >>
rect 145498 44513 145732 44519
rect 145498 44423 145505 44513
rect 145725 44423 145732 44513
rect 136996 44211 137230 44214
rect 136996 43983 136999 44211
rect 137227 43983 137230 44211
rect 136996 43911 137230 43983
rect 145498 44211 145732 44423
rect 145498 43983 145501 44211
rect 145729 43983 145732 44211
rect 145498 43375 145732 43983
rect 136996 38782 137230 38923
rect 139682 38814 142402 43375
rect 139682 38770 139916 38814
rect 145498 37591 145732 38932
rect 144959 37586 145732 37591
rect 144959 37362 144964 37586
rect 145150 37362 145732 37586
rect 144959 37357 145732 37362
rect 136164 35602 136398 35607
rect 136164 35379 136169 35602
rect 136392 35379 136398 35602
rect 136164 34705 136398 35379
rect 136996 35601 137230 36198
rect 136996 35378 137002 35601
rect 137225 35378 137230 35601
rect 138058 35681 138699 36145
rect 138058 35430 138102 35681
rect 138671 35430 138699 35681
rect 138058 35425 138699 35430
rect 136996 35373 137230 35378
rect 136164 34615 136171 34705
rect 136391 34615 136398 34705
rect 136164 34612 136398 34615
rect 136164 25214 136398 25218
rect 136164 25124 136171 25214
rect 136391 25124 136398 25214
rect 136164 23397 136398 25124
rect 138046 24669 138687 24683
rect 138046 24418 138090 24669
rect 138659 24418 138687 24669
rect 138046 23397 138687 24418
rect 136164 23207 136399 23397
rect 137171 23207 137177 23397
rect 136164 22951 137177 23207
rect 137171 22756 137177 22951
rect 138280 22756 138687 23397
rect 149309 23739 149703 23838
rect 149309 23249 149354 23739
rect 149698 23249 149703 23739
rect 149309 23216 149703 23249
rect 149684 23155 149703 23216
rect 139304 22923 139709 22928
rect 139304 22433 139309 22923
rect 139704 22433 139709 22923
rect 139304 22428 139709 22433
<< via2 >>
rect 145505 44423 145725 44513
rect 144964 37362 145150 37586
rect 138102 35430 138671 35681
rect 136171 34615 136391 34705
rect 136171 25124 136391 25214
rect 138090 24418 138659 24669
rect 149354 23249 149355 23739
rect 149355 23249 149697 23739
rect 139309 22433 139704 22923
<< metal3 >>
rect 145498 44513 145732 44519
rect 145498 44423 145505 44513
rect 145725 44423 145732 44513
rect 145498 44420 145732 44423
rect 144959 37586 145155 37591
rect 144959 37362 144964 37586
rect 145150 37362 145155 37586
rect 144959 37357 145155 37362
rect 138094 35681 138678 35686
rect 138094 35430 138102 35681
rect 138671 35430 138678 35681
rect 138094 35425 138678 35430
rect 136164 34705 136398 34709
rect 136164 34615 136171 34705
rect 136391 34615 136398 34705
rect 136164 34612 136398 34615
rect 136164 25214 136398 25218
rect 136164 25124 136171 25214
rect 136391 25124 136398 25214
rect 136164 25121 136398 25124
rect 138082 24669 138666 24674
rect 138082 24418 138090 24669
rect 138659 24418 138666 24669
rect 138082 24413 138666 24418
rect 149309 23739 149703 23838
rect 149309 23249 149354 23739
rect 149697 23249 149703 23739
rect 149309 23216 149703 23249
rect 139304 22923 139709 22928
rect 139304 22433 139309 22923
rect 139704 22433 139709 22923
rect 139304 22428 139709 22433
<< via3 >>
rect 145505 44423 145725 44513
rect 144964 37362 145150 37586
rect 138102 35430 138671 35681
rect 136171 34615 136391 34705
rect 136171 25124 136391 25214
rect 138090 24418 138659 24669
rect 149354 23249 149697 23739
rect 139309 22433 139704 22923
<< metal4 >>
rect 142409 54139 148798 54424
rect 142409 51123 145346 54139
rect 142409 44601 145369 51123
rect 145498 44513 145732 53916
rect 145861 51123 148798 54139
rect 145861 44602 148821 51123
rect 145498 44423 145505 44513
rect 145725 44423 145732 44513
rect 145498 44420 145732 44423
rect 144959 37586 145155 37591
rect 144959 37362 144964 37586
rect 145150 37362 145155 37586
rect 144959 37142 145155 37362
rect 138058 35681 138699 35688
rect 138058 35430 138102 35681
rect 138671 35430 138699 35681
rect 138058 35120 138699 35430
rect 133075 34835 139464 35120
rect 133075 31819 136012 34835
rect 136164 34705 136398 34709
rect 136164 34615 136171 34705
rect 136391 34615 136398 34705
rect 133075 25297 136035 31819
rect 136164 25214 136398 34615
rect 136527 31819 139464 34835
rect 140109 33443 140169 33943
rect 136527 30156 139487 31819
rect 136527 29798 139507 30156
rect 136527 25298 139487 29798
rect 136164 25124 136171 25214
rect 136391 25124 136398 25214
rect 136164 25121 136398 25124
rect 138046 24669 138687 25298
rect 138046 24418 138090 24669
rect 138659 24418 138687 24669
rect 138046 24411 138687 24418
rect 149350 23838 149703 23894
rect 149309 23739 149703 23838
rect 149309 23249 149354 23739
rect 149697 23249 149703 23739
rect 149309 23154 149703 23249
rect 149350 23149 149703 23154
rect 139304 22923 140139 22928
rect 139304 22433 139309 22923
rect 139704 22433 140139 22923
rect 139304 22428 140139 22433
use load_modulation  load_modulation_0
timestamp 1681069304
transform 0 1 137207 -1 0 23184
box -213 -36 428 1073
use rectifier  rectifier_0
timestamp 1681339707
transform 0 -1 148298 1 0 20477
box -2621 -1052 18329 8189
use resonator  resonator_0
timestamp 1682034855
transform 1 0 587701 0 1 -32688
box -586971 27283 -298971 375283
use ring_oscillator  ring_oscillator_0
timestamp 1681575212
transform 0 1 139571 -1 0 39555
box 755 -2575 3401 345
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_0
timestamp 1682220957
transform 1 0 134628 0 1 26778
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_1
timestamp 1682220957
transform 1 0 134628 0 1 29938
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_2
timestamp 1682220957
transform -1 0 137934 0 1 26778
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_3
timestamp 1682220957
transform -1 0 137934 0 1 29938
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_4
timestamp 1682220957
transform 1 0 134628 0 1 33098
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_5
timestamp 1682220957
transform -1 0 137934 0 1 33098
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_6
timestamp 1682220957
transform 1 0 143962 0 1 52402
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_7
timestamp 1682220957
transform -1 0 147268 0 1 52402
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_8
timestamp 1682220957
transform 1 0 143962 0 1 46082
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_9
timestamp 1682220957
transform 1 0 143962 0 1 49242
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_10
timestamp 1682220957
transform -1 0 147268 0 1 46082
box -1593 -1520 1593 1520
use sky130_fd_pr__cap_mim_m3_1_LJ5JLG  sky130_fd_pr__cap_mim_m3_1_LJ5JLG_11
timestamp 1682220957
transform -1 0 147268 0 1 49242
box -1593 -1520 1593 1520
use Temperature_Sensor  Temperature_Sensor_0
timestamp 1682114810
transform 0 1 139884 -1 0 40988
box -2924 -2888 2174 32
use voltage_limiter  voltage_limiter_0
timestamp 1682257554
transform 0 -1 141941 1 0 38473
box 329 -3791 4902 -446
<< end >>
