magic
tech sky130A
magscale 1 2
timestamp 1681382244
<< nwell >>
rect -294 -564 294 598
<< pmoslvt >>
rect -200 -464 200 536
<< pdiff >>
rect -258 524 -200 536
rect -258 -452 -246 524
rect -212 -452 -200 524
rect -258 -464 -200 -452
rect 200 524 258 536
rect 200 -452 212 524
rect 246 -452 258 524
rect 200 -464 258 -452
<< pdiffc >>
rect -246 -452 -212 524
rect 212 -452 246 524
<< poly >>
rect -200 536 200 562
rect -200 -511 200 -464
rect -200 -545 -184 -511
rect 184 -545 200 -511
rect -200 -561 200 -545
<< polycont >>
rect -184 -545 184 -511
<< locali >>
rect -246 524 -212 540
rect -246 -468 -212 -452
rect 212 524 246 540
rect 212 -468 246 -452
rect -200 -545 -184 -511
rect 184 -545 200 -511
<< viali >>
rect -246 -452 -212 524
rect 212 -452 246 524
rect -184 -545 184 -511
<< metal1 >>
rect -252 524 -206 536
rect -252 -452 -246 524
rect -212 -452 -206 524
rect -252 -464 -206 -452
rect 206 524 252 536
rect 206 -452 212 524
rect 246 -452 252 524
rect 206 -464 252 -452
rect -196 -511 196 -505
rect -196 -545 -184 -511
rect 184 -545 196 -511
rect -196 -551 196 -545
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
