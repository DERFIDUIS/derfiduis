** sch_path: /home/karlajcm/Documentos/TESIS DE
*+ GRADO/WORK_IN_PROGRESS/My_xschem/voltage_limiter_tb.sch
**.subckt voltage_limiter_tb vdd vrec
*.iopin vdd
*.iopin vrec
V1 vrec GND 1.8
.save i(v1)
x1 vrec GND vdd voltage_limiter


**** begin user architecture code

.control
save all
dc V1 0 3 0.01
plot vdd
set wr_singlescale
set wr_vecnames
wrdata vl_ll.txt v(vdd)
.endc


** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice ll


**** end user architecture code
**.ends

.include voltage_limiter.spice

.GLOBAL GND
.end
