magic
tech sky130A
magscale 1 2
timestamp 1681226341
<< nmoslvt >>
rect -200 -231 200 169
<< ndiff >>
rect -258 157 -200 169
rect -258 -219 -246 157
rect -212 -219 -200 157
rect -258 -231 -200 -219
rect 200 157 258 169
rect 200 -219 212 157
rect 246 -219 258 157
rect 200 -231 258 -219
<< ndiffc >>
rect -246 -219 -212 157
rect 212 -219 246 157
<< poly >>
rect -200 241 200 257
rect -200 207 -184 241
rect 184 207 200 241
rect -200 169 200 207
rect -200 -257 200 -231
<< polycont >>
rect -184 207 184 241
<< locali >>
rect -200 207 -184 241
rect 184 207 200 241
rect -246 157 -212 173
rect -246 -235 -212 -219
rect 212 157 246 173
rect 212 -235 246 -219
<< viali >>
rect -184 207 184 241
rect -246 -219 -212 157
rect 212 -219 246 157
<< metal1 >>
rect -196 241 196 247
rect -196 207 -184 241
rect 184 207 196 241
rect -196 201 196 207
rect -252 157 -206 169
rect -252 -219 -246 157
rect -212 -219 -206 157
rect -252 -231 -206 -219
rect 206 157 252 169
rect 206 -219 212 157
rect 246 -219 252 157
rect 206 -231 252 -219
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
