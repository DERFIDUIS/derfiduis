magic
tech sky130A
magscale 1 2
timestamp 1681224397
<< error_p >>
rect -294 -598 294 564
<< nwell >>
rect -294 -598 294 564
<< pmoslvt >>
rect -200 -536 200 464
<< pdiff >>
rect -258 452 -200 464
rect -258 -524 -246 452
rect -212 -524 -200 452
rect -258 -536 -200 -524
rect 200 452 258 464
rect 200 -524 212 452
rect 246 -524 258 452
rect 200 -536 258 -524
<< pdiffc >>
rect -246 -524 -212 452
rect 212 -524 246 452
<< poly >>
rect -200 545 200 561
rect -200 511 -184 545
rect 184 511 200 545
rect -200 464 200 511
rect -200 -562 200 -536
<< polycont >>
rect -184 511 184 545
<< locali >>
rect -200 511 -184 545
rect 184 511 200 545
rect -246 452 -212 468
rect -246 -540 -212 -524
rect 212 452 246 468
rect 212 -540 246 -524
<< viali >>
rect -184 511 184 545
rect -246 -524 -212 452
rect 212 -524 246 452
<< metal1 >>
rect -196 545 196 551
rect -196 511 -184 545
rect 184 511 196 545
rect -196 505 196 511
rect -252 452 -206 464
rect -252 -524 -246 452
rect -212 -524 -206 452
rect -252 -536 -206 -524
rect 206 452 252 464
rect 206 -524 212 452
rect 246 -524 252 452
rect 206 -536 252 -524
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
