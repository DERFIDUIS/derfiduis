magic
tech sky130A
magscale 1 2
timestamp 1680390383
<< xpolycontact >>
rect -141 282 141 714
rect -141 -714 141 -282
<< xpolyres >>
rect -141 -282 141 282
<< viali >>
rect -125 299 125 696
rect -125 -696 125 -299
<< metal1 >>
rect -131 696 131 708
rect -131 299 -125 696
rect 125 299 131 696
rect -131 287 131 299
rect -131 -299 131 -287
rect -131 -696 -125 -299
rect 125 -696 131 -299
rect -131 -708 131 -696
<< res1p41 >>
rect -143 -284 143 284
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 2.82 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 4.266k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
