magic
tech sky130A
magscale 1 2
timestamp 1681965435
<< nwell >>
rect 5168 -1712 5686 -1674
rect 3568 -2674 3634 -1712
rect 3976 -2674 4086 -1712
rect 4570 -1734 4682 -1712
rect 4570 -2674 4698 -1734
rect 5168 -1766 5234 -1712
rect 5620 -1766 5686 -1712
rect 5168 -1918 5686 -1766
rect 5168 -1956 5456 -1918
rect 5168 -2674 5234 -1956
rect 5620 -2674 5686 -1918
rect 6160 -2674 6284 -1712
rect 6768 -2674 6882 -1712
rect 7220 -2674 7286 -1712
<< pwell >>
rect 2358 -4610 2582 -1454
rect 2648 -6808 2882 -3124
rect 3250 -6808 3482 -3124
rect 3852 -6808 4086 -3124
rect 4454 -3586 4704 -3124
rect 4454 -6808 4688 -3586
rect 6010 -6808 6242 -3124
rect 6614 -6808 6848 -3124
rect 7218 -6808 7452 -3124
rect 7822 -6808 8058 -3124
rect 8426 -6808 8660 -3124
rect 9030 -6808 9262 -3124
<< ndiff >>
rect 5554 -5094 5556 -4694
<< pdiff >>
rect 3668 -2612 3670 -1812
rect 3984 -2612 3986 -1812
rect 4072 -2612 4074 -1812
rect 4690 -2612 4692 -1812
rect 5268 -2612 5270 -1812
rect 5584 -2612 5586 -1812
rect 6162 -2612 6164 -1812
rect 6780 -2612 6782 -1812
rect 6868 -2612 6870 -1812
rect 7184 -2612 7186 -1812
<< psubdiff >>
rect 2454 -1616 2582 -1454
rect 2454 -1788 2478 -1616
rect 2558 -1788 2582 -1616
rect 2454 -1888 2582 -1788
rect 2454 -2060 2478 -1888
rect 2558 -2060 2582 -1888
rect 2454 -2222 2582 -2060
rect 2454 -2394 2478 -2222
rect 2558 -2394 2582 -2222
rect 2454 -2534 2582 -2394
rect 2454 -2706 2478 -2534
rect 2558 -2706 2582 -2534
rect 2454 -2840 2582 -2706
rect 2454 -3012 2478 -2840
rect 2558 -3012 2582 -2840
rect 2454 -3098 2582 -3012
rect 2454 -3270 2478 -3098
rect 2558 -3270 2582 -3098
rect 2454 -3370 2582 -3270
rect 2454 -3542 2478 -3370
rect 2558 -3542 2582 -3370
rect 2454 -3704 2582 -3542
rect 2454 -3876 2478 -3704
rect 2558 -3876 2582 -3704
rect 2454 -4016 2582 -3876
rect 2454 -4188 2478 -4016
rect 2558 -4188 2582 -4016
rect 2454 -4322 2582 -4188
rect 2454 -4494 2478 -4322
rect 2558 -4494 2582 -4322
rect 2454 -4610 2582 -4494
rect 2648 -3240 2776 -3124
rect 2648 -3412 2672 -3240
rect 2752 -3412 2776 -3240
rect 2648 -3512 2776 -3412
rect 2648 -3684 2672 -3512
rect 2752 -3684 2776 -3512
rect 2648 -3822 2776 -3684
rect 2648 -3994 2672 -3822
rect 2752 -3994 2776 -3822
rect 2648 -4094 2776 -3994
rect 2648 -4266 2672 -4094
rect 2752 -4266 2776 -4094
rect 2648 -4428 2776 -4266
rect 2648 -4600 2672 -4428
rect 2752 -4600 2776 -4428
rect 2648 -4740 2776 -4600
rect 2648 -4912 2672 -4740
rect 2752 -4912 2776 -4740
rect 2648 -5046 2776 -4912
rect 2648 -5218 2672 -5046
rect 2752 -5218 2776 -5046
rect 2648 -5332 2776 -5218
rect 2648 -5504 2672 -5332
rect 2752 -5504 2776 -5332
rect 2648 -5604 2776 -5504
rect 2648 -5776 2672 -5604
rect 2752 -5776 2776 -5604
rect 2648 -5938 2776 -5776
rect 2648 -6110 2672 -5938
rect 2752 -6110 2776 -5938
rect 2648 -6250 2776 -6110
rect 2648 -6422 2672 -6250
rect 2752 -6422 2776 -6250
rect 2648 -6556 2776 -6422
rect 2648 -6728 2672 -6556
rect 2752 -6728 2776 -6556
rect 2648 -6808 2776 -6728
rect 3250 -3240 3378 -3124
rect 3250 -3412 3274 -3240
rect 3354 -3412 3378 -3240
rect 3250 -3512 3378 -3412
rect 3250 -3684 3274 -3512
rect 3354 -3684 3378 -3512
rect 3250 -3822 3378 -3684
rect 3250 -3994 3274 -3822
rect 3354 -3994 3378 -3822
rect 3250 -4094 3378 -3994
rect 3250 -4266 3274 -4094
rect 3354 -4266 3378 -4094
rect 3250 -4428 3378 -4266
rect 3250 -4600 3274 -4428
rect 3354 -4600 3378 -4428
rect 3250 -4740 3378 -4600
rect 3250 -4912 3274 -4740
rect 3354 -4912 3378 -4740
rect 3250 -5046 3378 -4912
rect 3250 -5218 3274 -5046
rect 3354 -5218 3378 -5046
rect 3250 -5332 3378 -5218
rect 3250 -5504 3274 -5332
rect 3354 -5504 3378 -5332
rect 3250 -5604 3378 -5504
rect 3250 -5776 3274 -5604
rect 3354 -5776 3378 -5604
rect 3250 -5938 3378 -5776
rect 3250 -6110 3274 -5938
rect 3354 -6110 3378 -5938
rect 3250 -6250 3378 -6110
rect 3250 -6422 3274 -6250
rect 3354 -6422 3378 -6250
rect 3250 -6556 3378 -6422
rect 3250 -6728 3274 -6556
rect 3354 -6728 3378 -6556
rect 3250 -6808 3378 -6728
rect 3852 -3240 3980 -3124
rect 3852 -3412 3876 -3240
rect 3956 -3412 3980 -3240
rect 3852 -3512 3980 -3412
rect 3852 -3684 3876 -3512
rect 3956 -3684 3980 -3512
rect 3852 -3822 3980 -3684
rect 3852 -3994 3876 -3822
rect 3956 -3994 3980 -3822
rect 3852 -4094 3980 -3994
rect 3852 -4266 3876 -4094
rect 3956 -4266 3980 -4094
rect 3852 -4428 3980 -4266
rect 3852 -4600 3876 -4428
rect 3956 -4600 3980 -4428
rect 3852 -4740 3980 -4600
rect 3852 -4912 3876 -4740
rect 3956 -4912 3980 -4740
rect 3852 -5046 3980 -4912
rect 3852 -5218 3876 -5046
rect 3956 -5218 3980 -5046
rect 3852 -5332 3980 -5218
rect 3852 -5504 3876 -5332
rect 3956 -5504 3980 -5332
rect 3852 -5604 3980 -5504
rect 3852 -5776 3876 -5604
rect 3956 -5776 3980 -5604
rect 3852 -5938 3980 -5776
rect 3852 -6110 3876 -5938
rect 3956 -6110 3980 -5938
rect 3852 -6250 3980 -6110
rect 3852 -6422 3876 -6250
rect 3956 -6422 3980 -6250
rect 3852 -6556 3980 -6422
rect 3852 -6728 3876 -6556
rect 3956 -6728 3980 -6556
rect 3852 -6808 3980 -6728
rect 4454 -3240 4582 -3124
rect 4454 -3412 4478 -3240
rect 4558 -3412 4582 -3240
rect 4454 -3512 4582 -3412
rect 4454 -3684 4478 -3512
rect 4558 -3684 4582 -3512
rect 4454 -3822 4582 -3684
rect 4454 -3994 4478 -3822
rect 4558 -3994 4582 -3822
rect 4454 -4094 4582 -3994
rect 4454 -4266 4478 -4094
rect 4558 -4266 4582 -4094
rect 4454 -4428 4582 -4266
rect 4454 -4600 4478 -4428
rect 4558 -4600 4582 -4428
rect 4454 -4740 4582 -4600
rect 6010 -3240 6138 -3124
rect 6010 -3412 6034 -3240
rect 6114 -3412 6138 -3240
rect 6010 -3512 6138 -3412
rect 6010 -3684 6034 -3512
rect 6114 -3684 6138 -3512
rect 6010 -3822 6138 -3684
rect 6010 -3994 6034 -3822
rect 6114 -3994 6138 -3822
rect 6010 -4094 6138 -3994
rect 6010 -4266 6034 -4094
rect 6114 -4266 6138 -4094
rect 6010 -4428 6138 -4266
rect 6010 -4600 6034 -4428
rect 6114 -4600 6138 -4428
rect 4454 -4912 4478 -4740
rect 4558 -4912 4582 -4740
rect 4454 -5046 4582 -4912
rect 4454 -5218 4478 -5046
rect 4558 -5218 4582 -5046
rect 5556 -4760 5620 -4694
rect 5556 -4794 5582 -4760
rect 5616 -4794 5620 -4760
rect 5556 -4828 5620 -4794
rect 5556 -4862 5582 -4828
rect 5616 -4862 5620 -4828
rect 5556 -4896 5620 -4862
rect 5556 -4930 5582 -4896
rect 5616 -4930 5620 -4896
rect 5556 -4964 5620 -4930
rect 5556 -4998 5582 -4964
rect 5616 -4998 5620 -4964
rect 5556 -5032 5620 -4998
rect 5556 -5066 5582 -5032
rect 5616 -5066 5620 -5032
rect 5556 -5094 5620 -5066
rect 6010 -4740 6138 -4600
rect 6010 -4912 6034 -4740
rect 6114 -4912 6138 -4740
rect 6010 -5046 6138 -4912
rect 4454 -5332 4582 -5218
rect 4454 -5504 4478 -5332
rect 4558 -5504 4582 -5332
rect 4454 -5604 4582 -5504
rect 4454 -5776 4478 -5604
rect 4558 -5776 4582 -5604
rect 4454 -5938 4582 -5776
rect 4454 -6110 4478 -5938
rect 4558 -6110 4582 -5938
rect 4454 -6250 4582 -6110
rect 4454 -6422 4478 -6250
rect 4558 -6422 4582 -6250
rect 4454 -6556 4582 -6422
rect 4454 -6728 4478 -6556
rect 4558 -6728 4582 -6556
rect 4454 -6808 4582 -6728
rect 6010 -5218 6034 -5046
rect 6114 -5218 6138 -5046
rect 6010 -5332 6138 -5218
rect 6010 -5504 6034 -5332
rect 6114 -5504 6138 -5332
rect 6010 -5604 6138 -5504
rect 6010 -5776 6034 -5604
rect 6114 -5776 6138 -5604
rect 6010 -5938 6138 -5776
rect 6010 -6110 6034 -5938
rect 6114 -6110 6138 -5938
rect 6010 -6250 6138 -6110
rect 6010 -6422 6034 -6250
rect 6114 -6422 6138 -6250
rect 6010 -6556 6138 -6422
rect 6010 -6728 6034 -6556
rect 6114 -6728 6138 -6556
rect 6010 -6808 6138 -6728
rect 6614 -3240 6742 -3124
rect 6614 -3412 6638 -3240
rect 6718 -3412 6742 -3240
rect 6614 -3512 6742 -3412
rect 6614 -3684 6638 -3512
rect 6718 -3684 6742 -3512
rect 6614 -3822 6742 -3684
rect 6614 -3994 6638 -3822
rect 6718 -3994 6742 -3822
rect 6614 -4094 6742 -3994
rect 6614 -4266 6638 -4094
rect 6718 -4266 6742 -4094
rect 6614 -4428 6742 -4266
rect 6614 -4600 6638 -4428
rect 6718 -4600 6742 -4428
rect 6614 -4740 6742 -4600
rect 6614 -4912 6638 -4740
rect 6718 -4912 6742 -4740
rect 6614 -5046 6742 -4912
rect 6614 -5218 6638 -5046
rect 6718 -5218 6742 -5046
rect 6614 -5332 6742 -5218
rect 6614 -5504 6638 -5332
rect 6718 -5504 6742 -5332
rect 6614 -5604 6742 -5504
rect 6614 -5776 6638 -5604
rect 6718 -5776 6742 -5604
rect 6614 -5938 6742 -5776
rect 6614 -6110 6638 -5938
rect 6718 -6110 6742 -5938
rect 6614 -6250 6742 -6110
rect 6614 -6422 6638 -6250
rect 6718 -6422 6742 -6250
rect 6614 -6556 6742 -6422
rect 6614 -6728 6638 -6556
rect 6718 -6728 6742 -6556
rect 6614 -6808 6742 -6728
rect 7218 -3240 7346 -3124
rect 7218 -3412 7242 -3240
rect 7322 -3412 7346 -3240
rect 7218 -3512 7346 -3412
rect 7218 -3684 7242 -3512
rect 7322 -3684 7346 -3512
rect 7218 -3822 7346 -3684
rect 7218 -3994 7242 -3822
rect 7322 -3994 7346 -3822
rect 7218 -4094 7346 -3994
rect 7218 -4266 7242 -4094
rect 7322 -4266 7346 -4094
rect 7218 -4428 7346 -4266
rect 7218 -4600 7242 -4428
rect 7322 -4600 7346 -4428
rect 7218 -4740 7346 -4600
rect 7218 -4912 7242 -4740
rect 7322 -4912 7346 -4740
rect 7218 -5046 7346 -4912
rect 7218 -5218 7242 -5046
rect 7322 -5218 7346 -5046
rect 7218 -5332 7346 -5218
rect 7218 -5504 7242 -5332
rect 7322 -5504 7346 -5332
rect 7218 -5604 7346 -5504
rect 7218 -5776 7242 -5604
rect 7322 -5776 7346 -5604
rect 7218 -5938 7346 -5776
rect 7218 -6110 7242 -5938
rect 7322 -6110 7346 -5938
rect 7218 -6250 7346 -6110
rect 7218 -6422 7242 -6250
rect 7322 -6422 7346 -6250
rect 7218 -6556 7346 -6422
rect 7218 -6728 7242 -6556
rect 7322 -6728 7346 -6556
rect 7218 -6808 7346 -6728
rect 7822 -3240 7950 -3124
rect 7822 -3412 7846 -3240
rect 7926 -3412 7950 -3240
rect 7822 -3512 7950 -3412
rect 7822 -3684 7846 -3512
rect 7926 -3684 7950 -3512
rect 7822 -3822 7950 -3684
rect 7822 -3994 7846 -3822
rect 7926 -3994 7950 -3822
rect 7822 -4094 7950 -3994
rect 7822 -4266 7846 -4094
rect 7926 -4266 7950 -4094
rect 7822 -4428 7950 -4266
rect 7822 -4600 7846 -4428
rect 7926 -4600 7950 -4428
rect 7822 -4740 7950 -4600
rect 7822 -4912 7846 -4740
rect 7926 -4912 7950 -4740
rect 7822 -5046 7950 -4912
rect 7822 -5218 7846 -5046
rect 7926 -5218 7950 -5046
rect 7822 -5332 7950 -5218
rect 7822 -5504 7846 -5332
rect 7926 -5504 7950 -5332
rect 7822 -5604 7950 -5504
rect 7822 -5776 7846 -5604
rect 7926 -5776 7950 -5604
rect 7822 -5938 7950 -5776
rect 7822 -6110 7846 -5938
rect 7926 -6110 7950 -5938
rect 7822 -6250 7950 -6110
rect 7822 -6422 7846 -6250
rect 7926 -6422 7950 -6250
rect 7822 -6556 7950 -6422
rect 7822 -6728 7846 -6556
rect 7926 -6728 7950 -6556
rect 7822 -6808 7950 -6728
rect 8426 -3240 8554 -3124
rect 8426 -3412 8450 -3240
rect 8530 -3412 8554 -3240
rect 8426 -3512 8554 -3412
rect 8426 -3684 8450 -3512
rect 8530 -3684 8554 -3512
rect 8426 -3822 8554 -3684
rect 8426 -3994 8450 -3822
rect 8530 -3994 8554 -3822
rect 8426 -4094 8554 -3994
rect 8426 -4266 8450 -4094
rect 8530 -4266 8554 -4094
rect 8426 -4428 8554 -4266
rect 8426 -4600 8450 -4428
rect 8530 -4600 8554 -4428
rect 8426 -4740 8554 -4600
rect 8426 -4912 8450 -4740
rect 8530 -4912 8554 -4740
rect 8426 -5046 8554 -4912
rect 8426 -5218 8450 -5046
rect 8530 -5218 8554 -5046
rect 8426 -5332 8554 -5218
rect 8426 -5504 8450 -5332
rect 8530 -5504 8554 -5332
rect 8426 -5604 8554 -5504
rect 8426 -5776 8450 -5604
rect 8530 -5776 8554 -5604
rect 8426 -5938 8554 -5776
rect 8426 -6110 8450 -5938
rect 8530 -6110 8554 -5938
rect 8426 -6250 8554 -6110
rect 8426 -6422 8450 -6250
rect 8530 -6422 8554 -6250
rect 8426 -6556 8554 -6422
rect 8426 -6728 8450 -6556
rect 8530 -6728 8554 -6556
rect 8426 -6808 8554 -6728
rect 9030 -3240 9158 -3124
rect 9030 -3412 9054 -3240
rect 9134 -3412 9158 -3240
rect 9030 -3512 9158 -3412
rect 9030 -3684 9054 -3512
rect 9134 -3684 9158 -3512
rect 9030 -3822 9158 -3684
rect 9030 -3994 9054 -3822
rect 9134 -3994 9158 -3822
rect 9030 -4094 9158 -3994
rect 9030 -4266 9054 -4094
rect 9134 -4266 9158 -4094
rect 9030 -4428 9158 -4266
rect 9030 -4600 9054 -4428
rect 9134 -4600 9158 -4428
rect 9030 -4740 9158 -4600
rect 9030 -4912 9054 -4740
rect 9134 -4912 9158 -4740
rect 9030 -5046 9158 -4912
rect 9030 -5218 9054 -5046
rect 9134 -5218 9158 -5046
rect 9030 -5332 9158 -5218
rect 9030 -5504 9054 -5332
rect 9134 -5504 9158 -5332
rect 9030 -5604 9158 -5504
rect 9030 -5776 9054 -5604
rect 9134 -5776 9158 -5604
rect 9030 -5938 9158 -5776
rect 9030 -6110 9054 -5938
rect 9134 -6110 9158 -5938
rect 9030 -6250 9158 -6110
rect 9030 -6422 9054 -6250
rect 9134 -6422 9158 -6250
rect 9030 -6556 9158 -6422
rect 9030 -6728 9054 -6556
rect 9134 -6728 9158 -6556
rect 9030 -6808 9158 -6728
<< nsubdiff >>
rect 3604 -1840 3668 -1812
rect 3604 -1874 3608 -1840
rect 3642 -1874 3668 -1840
rect 3604 -1908 3668 -1874
rect 3604 -1942 3608 -1908
rect 3642 -1942 3668 -1908
rect 3604 -1976 3668 -1942
rect 3604 -2010 3608 -1976
rect 3642 -2010 3668 -1976
rect 3604 -2044 3668 -2010
rect 3604 -2078 3608 -2044
rect 3642 -2078 3668 -2044
rect 3604 -2112 3668 -2078
rect 3604 -2146 3608 -2112
rect 3642 -2146 3668 -2112
rect 3604 -2180 3668 -2146
rect 3604 -2214 3608 -2180
rect 3642 -2214 3668 -2180
rect 3604 -2248 3668 -2214
rect 3604 -2282 3608 -2248
rect 3642 -2282 3668 -2248
rect 3604 -2316 3668 -2282
rect 3604 -2350 3608 -2316
rect 3642 -2350 3668 -2316
rect 3604 -2384 3668 -2350
rect 3604 -2418 3608 -2384
rect 3642 -2418 3668 -2384
rect 3604 -2452 3668 -2418
rect 3604 -2486 3608 -2452
rect 3642 -2486 3668 -2452
rect 3604 -2520 3668 -2486
rect 3604 -2554 3608 -2520
rect 3642 -2554 3668 -2520
rect 3604 -2612 3668 -2554
rect 3986 -1840 4072 -1812
rect 3986 -1874 4012 -1840
rect 4046 -1874 4072 -1840
rect 3986 -1908 4072 -1874
rect 3986 -1942 4012 -1908
rect 4046 -1942 4072 -1908
rect 3986 -1976 4072 -1942
rect 3986 -2010 4012 -1976
rect 4046 -2010 4072 -1976
rect 3986 -2044 4072 -2010
rect 3986 -2078 4012 -2044
rect 4046 -2078 4072 -2044
rect 3986 -2112 4072 -2078
rect 3986 -2146 4012 -2112
rect 4046 -2146 4072 -2112
rect 3986 -2180 4072 -2146
rect 3986 -2214 4012 -2180
rect 4046 -2214 4072 -2180
rect 3986 -2248 4072 -2214
rect 3986 -2282 4012 -2248
rect 4046 -2282 4072 -2248
rect 3986 -2316 4072 -2282
rect 3986 -2350 4012 -2316
rect 4046 -2350 4072 -2316
rect 3986 -2384 4072 -2350
rect 3986 -2418 4012 -2384
rect 4046 -2418 4072 -2384
rect 3986 -2452 4072 -2418
rect 3986 -2486 4012 -2452
rect 4046 -2486 4072 -2452
rect 3986 -2520 4072 -2486
rect 3986 -2554 4012 -2520
rect 4046 -2554 4072 -2520
rect 3986 -2612 4072 -2554
rect 4606 -1840 4690 -1812
rect 4606 -1874 4610 -1840
rect 4644 -1874 4690 -1840
rect 4606 -1908 4690 -1874
rect 4606 -1942 4610 -1908
rect 4644 -1942 4690 -1908
rect 4606 -1976 4690 -1942
rect 4606 -2010 4610 -1976
rect 4644 -2010 4690 -1976
rect 4606 -2044 4690 -2010
rect 4606 -2078 4610 -2044
rect 4644 -2078 4690 -2044
rect 4606 -2112 4690 -2078
rect 4606 -2146 4610 -2112
rect 4644 -2146 4690 -2112
rect 4606 -2180 4690 -2146
rect 4606 -2214 4610 -2180
rect 4644 -2214 4690 -2180
rect 4606 -2248 4690 -2214
rect 4606 -2282 4610 -2248
rect 4644 -2282 4690 -2248
rect 4606 -2316 4690 -2282
rect 4606 -2350 4610 -2316
rect 4644 -2350 4690 -2316
rect 4606 -2384 4690 -2350
rect 4606 -2418 4610 -2384
rect 4644 -2418 4690 -2384
rect 4606 -2452 4690 -2418
rect 4606 -2486 4610 -2452
rect 4644 -2486 4690 -2452
rect 4606 -2520 4690 -2486
rect 4606 -2554 4610 -2520
rect 4644 -2554 4690 -2520
rect 4606 -2612 4690 -2554
rect 5204 -1870 5268 -1812
rect 5204 -1904 5208 -1870
rect 5242 -1904 5268 -1870
rect 5204 -1938 5268 -1904
rect 5204 -1972 5208 -1938
rect 5242 -1972 5268 -1938
rect 5204 -2006 5268 -1972
rect 5204 -2040 5208 -2006
rect 5242 -2040 5268 -2006
rect 5204 -2074 5268 -2040
rect 5204 -2108 5208 -2074
rect 5242 -2108 5268 -2074
rect 5204 -2142 5268 -2108
rect 5204 -2176 5208 -2142
rect 5242 -2176 5268 -2142
rect 5204 -2210 5268 -2176
rect 5204 -2244 5208 -2210
rect 5242 -2244 5268 -2210
rect 5204 -2278 5268 -2244
rect 5204 -2312 5208 -2278
rect 5242 -2312 5268 -2278
rect 5204 -2346 5268 -2312
rect 5204 -2380 5208 -2346
rect 5242 -2380 5268 -2346
rect 5204 -2414 5268 -2380
rect 5204 -2448 5208 -2414
rect 5242 -2448 5268 -2414
rect 5204 -2482 5268 -2448
rect 5204 -2516 5208 -2482
rect 5242 -2516 5268 -2482
rect 5204 -2550 5268 -2516
rect 5204 -2584 5208 -2550
rect 5242 -2584 5268 -2550
rect 5204 -2612 5268 -2584
rect 5586 -1870 5650 -1812
rect 5586 -1904 5612 -1870
rect 5646 -1904 5650 -1870
rect 5586 -1938 5650 -1904
rect 5586 -1972 5612 -1938
rect 5646 -1972 5650 -1938
rect 5586 -2006 5650 -1972
rect 5586 -2040 5612 -2006
rect 5646 -2040 5650 -2006
rect 5586 -2074 5650 -2040
rect 5586 -2108 5612 -2074
rect 5646 -2108 5650 -2074
rect 5586 -2142 5650 -2108
rect 5586 -2176 5612 -2142
rect 5646 -2176 5650 -2142
rect 5586 -2210 5650 -2176
rect 5586 -2244 5612 -2210
rect 5646 -2244 5650 -2210
rect 5586 -2278 5650 -2244
rect 5586 -2312 5612 -2278
rect 5646 -2312 5650 -2278
rect 5586 -2346 5650 -2312
rect 5586 -2380 5612 -2346
rect 5646 -2380 5650 -2346
rect 5586 -2414 5650 -2380
rect 5586 -2448 5612 -2414
rect 5646 -2448 5650 -2414
rect 5586 -2482 5650 -2448
rect 5586 -2516 5612 -2482
rect 5646 -2516 5650 -2482
rect 5586 -2550 5650 -2516
rect 5586 -2584 5612 -2550
rect 5646 -2584 5650 -2550
rect 5586 -2612 5650 -2584
rect 6164 -1840 6248 -1812
rect 6164 -1874 6210 -1840
rect 6244 -1874 6248 -1840
rect 6164 -1908 6248 -1874
rect 6164 -1942 6210 -1908
rect 6244 -1942 6248 -1908
rect 6164 -1976 6248 -1942
rect 6164 -2010 6210 -1976
rect 6244 -2010 6248 -1976
rect 6164 -2044 6248 -2010
rect 6164 -2078 6210 -2044
rect 6244 -2078 6248 -2044
rect 6164 -2112 6248 -2078
rect 6164 -2146 6210 -2112
rect 6244 -2146 6248 -2112
rect 6164 -2180 6248 -2146
rect 6164 -2214 6210 -2180
rect 6244 -2214 6248 -2180
rect 6164 -2248 6248 -2214
rect 6164 -2282 6210 -2248
rect 6244 -2282 6248 -2248
rect 6164 -2316 6248 -2282
rect 6164 -2350 6210 -2316
rect 6244 -2350 6248 -2316
rect 6164 -2384 6248 -2350
rect 6164 -2418 6210 -2384
rect 6244 -2418 6248 -2384
rect 6164 -2452 6248 -2418
rect 6164 -2486 6210 -2452
rect 6244 -2486 6248 -2452
rect 6164 -2520 6248 -2486
rect 6164 -2554 6210 -2520
rect 6244 -2554 6248 -2520
rect 6164 -2612 6248 -2554
rect 6782 -1840 6868 -1812
rect 6782 -1874 6808 -1840
rect 6842 -1874 6868 -1840
rect 6782 -1908 6868 -1874
rect 6782 -1942 6808 -1908
rect 6842 -1942 6868 -1908
rect 6782 -1976 6868 -1942
rect 6782 -2010 6808 -1976
rect 6842 -2010 6868 -1976
rect 6782 -2044 6868 -2010
rect 6782 -2078 6808 -2044
rect 6842 -2078 6868 -2044
rect 6782 -2112 6868 -2078
rect 6782 -2146 6808 -2112
rect 6842 -2146 6868 -2112
rect 6782 -2180 6868 -2146
rect 6782 -2214 6808 -2180
rect 6842 -2214 6868 -2180
rect 6782 -2248 6868 -2214
rect 6782 -2282 6808 -2248
rect 6842 -2282 6868 -2248
rect 6782 -2316 6868 -2282
rect 6782 -2350 6808 -2316
rect 6842 -2350 6868 -2316
rect 6782 -2384 6868 -2350
rect 6782 -2418 6808 -2384
rect 6842 -2418 6868 -2384
rect 6782 -2452 6868 -2418
rect 6782 -2486 6808 -2452
rect 6842 -2486 6868 -2452
rect 6782 -2520 6868 -2486
rect 6782 -2554 6808 -2520
rect 6842 -2554 6868 -2520
rect 6782 -2612 6868 -2554
rect 7186 -1840 7250 -1812
rect 7186 -1874 7212 -1840
rect 7246 -1874 7250 -1840
rect 7186 -1908 7250 -1874
rect 7186 -1942 7212 -1908
rect 7246 -1942 7250 -1908
rect 7186 -1976 7250 -1942
rect 7186 -2010 7212 -1976
rect 7246 -2010 7250 -1976
rect 7186 -2044 7250 -2010
rect 7186 -2078 7212 -2044
rect 7246 -2078 7250 -2044
rect 7186 -2112 7250 -2078
rect 7186 -2146 7212 -2112
rect 7246 -2146 7250 -2112
rect 7186 -2180 7250 -2146
rect 7186 -2214 7212 -2180
rect 7246 -2214 7250 -2180
rect 7186 -2248 7250 -2214
rect 7186 -2282 7212 -2248
rect 7246 -2282 7250 -2248
rect 7186 -2316 7250 -2282
rect 7186 -2350 7212 -2316
rect 7246 -2350 7250 -2316
rect 7186 -2384 7250 -2350
rect 7186 -2418 7212 -2384
rect 7246 -2418 7250 -2384
rect 7186 -2452 7250 -2418
rect 7186 -2486 7212 -2452
rect 7246 -2486 7250 -2452
rect 7186 -2520 7250 -2486
rect 7186 -2554 7212 -2520
rect 7246 -2554 7250 -2520
rect 7186 -2612 7250 -2554
<< psubdiffcont >>
rect 2478 -1788 2558 -1616
rect 2478 -2060 2558 -1888
rect 2478 -2394 2558 -2222
rect 2478 -2706 2558 -2534
rect 2478 -3012 2558 -2840
rect 2478 -3270 2558 -3098
rect 2478 -3542 2558 -3370
rect 2478 -3876 2558 -3704
rect 2478 -4188 2558 -4016
rect 2478 -4494 2558 -4322
rect 2672 -3412 2752 -3240
rect 2672 -3684 2752 -3512
rect 2672 -3994 2752 -3822
rect 2672 -4266 2752 -4094
rect 2672 -4600 2752 -4428
rect 2672 -4912 2752 -4740
rect 2672 -5218 2752 -5046
rect 2672 -5504 2752 -5332
rect 2672 -5776 2752 -5604
rect 2672 -6110 2752 -5938
rect 2672 -6422 2752 -6250
rect 2672 -6728 2752 -6556
rect 3274 -3412 3354 -3240
rect 3274 -3684 3354 -3512
rect 3274 -3994 3354 -3822
rect 3274 -4266 3354 -4094
rect 3274 -4600 3354 -4428
rect 3274 -4912 3354 -4740
rect 3274 -5218 3354 -5046
rect 3274 -5504 3354 -5332
rect 3274 -5776 3354 -5604
rect 3274 -6110 3354 -5938
rect 3274 -6422 3354 -6250
rect 3274 -6728 3354 -6556
rect 3876 -3412 3956 -3240
rect 3876 -3684 3956 -3512
rect 3876 -3994 3956 -3822
rect 3876 -4266 3956 -4094
rect 3876 -4600 3956 -4428
rect 3876 -4912 3956 -4740
rect 3876 -5218 3956 -5046
rect 3876 -5504 3956 -5332
rect 3876 -5776 3956 -5604
rect 3876 -6110 3956 -5938
rect 3876 -6422 3956 -6250
rect 3876 -6728 3956 -6556
rect 4478 -3412 4558 -3240
rect 4478 -3684 4558 -3512
rect 4478 -3994 4558 -3822
rect 4478 -4266 4558 -4094
rect 4478 -4600 4558 -4428
rect 6034 -3412 6114 -3240
rect 6034 -3684 6114 -3512
rect 6034 -3994 6114 -3822
rect 6034 -4266 6114 -4094
rect 6034 -4600 6114 -4428
rect 4478 -4912 4558 -4740
rect 4478 -5218 4558 -5046
rect 5582 -4794 5616 -4760
rect 5582 -4862 5616 -4828
rect 5582 -4930 5616 -4896
rect 5582 -4998 5616 -4964
rect 5582 -5066 5616 -5032
rect 6034 -4912 6114 -4740
rect 4478 -5504 4558 -5332
rect 4478 -5776 4558 -5604
rect 4478 -6110 4558 -5938
rect 4478 -6422 4558 -6250
rect 4478 -6728 4558 -6556
rect 6034 -5218 6114 -5046
rect 6034 -5504 6114 -5332
rect 6034 -5776 6114 -5604
rect 6034 -6110 6114 -5938
rect 6034 -6422 6114 -6250
rect 6034 -6728 6114 -6556
rect 6638 -3412 6718 -3240
rect 6638 -3684 6718 -3512
rect 6638 -3994 6718 -3822
rect 6638 -4266 6718 -4094
rect 6638 -4600 6718 -4428
rect 6638 -4912 6718 -4740
rect 6638 -5218 6718 -5046
rect 6638 -5504 6718 -5332
rect 6638 -5776 6718 -5604
rect 6638 -6110 6718 -5938
rect 6638 -6422 6718 -6250
rect 6638 -6728 6718 -6556
rect 7242 -3412 7322 -3240
rect 7242 -3684 7322 -3512
rect 7242 -3994 7322 -3822
rect 7242 -4266 7322 -4094
rect 7242 -4600 7322 -4428
rect 7242 -4912 7322 -4740
rect 7242 -5218 7322 -5046
rect 7242 -5504 7322 -5332
rect 7242 -5776 7322 -5604
rect 7242 -6110 7322 -5938
rect 7242 -6422 7322 -6250
rect 7242 -6728 7322 -6556
rect 7846 -3412 7926 -3240
rect 7846 -3684 7926 -3512
rect 7846 -3994 7926 -3822
rect 7846 -4266 7926 -4094
rect 7846 -4600 7926 -4428
rect 7846 -4912 7926 -4740
rect 7846 -5218 7926 -5046
rect 7846 -5504 7926 -5332
rect 7846 -5776 7926 -5604
rect 7846 -6110 7926 -5938
rect 7846 -6422 7926 -6250
rect 7846 -6728 7926 -6556
rect 8450 -3412 8530 -3240
rect 8450 -3684 8530 -3512
rect 8450 -3994 8530 -3822
rect 8450 -4266 8530 -4094
rect 8450 -4600 8530 -4428
rect 8450 -4912 8530 -4740
rect 8450 -5218 8530 -5046
rect 8450 -5504 8530 -5332
rect 8450 -5776 8530 -5604
rect 8450 -6110 8530 -5938
rect 8450 -6422 8530 -6250
rect 8450 -6728 8530 -6556
rect 9054 -3412 9134 -3240
rect 9054 -3684 9134 -3512
rect 9054 -3994 9134 -3822
rect 9054 -4266 9134 -4094
rect 9054 -4600 9134 -4428
rect 9054 -4912 9134 -4740
rect 9054 -5218 9134 -5046
rect 9054 -5504 9134 -5332
rect 9054 -5776 9134 -5604
rect 9054 -6110 9134 -5938
rect 9054 -6422 9134 -6250
rect 9054 -6728 9134 -6556
<< nsubdiffcont >>
rect 3608 -1874 3642 -1840
rect 3608 -1942 3642 -1908
rect 3608 -2010 3642 -1976
rect 3608 -2078 3642 -2044
rect 3608 -2146 3642 -2112
rect 3608 -2214 3642 -2180
rect 3608 -2282 3642 -2248
rect 3608 -2350 3642 -2316
rect 3608 -2418 3642 -2384
rect 3608 -2486 3642 -2452
rect 3608 -2554 3642 -2520
rect 4012 -1874 4046 -1840
rect 4012 -1942 4046 -1908
rect 4012 -2010 4046 -1976
rect 4012 -2078 4046 -2044
rect 4012 -2146 4046 -2112
rect 4012 -2214 4046 -2180
rect 4012 -2282 4046 -2248
rect 4012 -2350 4046 -2316
rect 4012 -2418 4046 -2384
rect 4012 -2486 4046 -2452
rect 4012 -2554 4046 -2520
rect 4610 -1874 4644 -1840
rect 4610 -1942 4644 -1908
rect 4610 -2010 4644 -1976
rect 4610 -2078 4644 -2044
rect 4610 -2146 4644 -2112
rect 4610 -2214 4644 -2180
rect 4610 -2282 4644 -2248
rect 4610 -2350 4644 -2316
rect 4610 -2418 4644 -2384
rect 4610 -2486 4644 -2452
rect 4610 -2554 4644 -2520
rect 5208 -1904 5242 -1870
rect 5208 -1972 5242 -1938
rect 5208 -2040 5242 -2006
rect 5208 -2108 5242 -2074
rect 5208 -2176 5242 -2142
rect 5208 -2244 5242 -2210
rect 5208 -2312 5242 -2278
rect 5208 -2380 5242 -2346
rect 5208 -2448 5242 -2414
rect 5208 -2516 5242 -2482
rect 5208 -2584 5242 -2550
rect 5612 -1904 5646 -1870
rect 5612 -1972 5646 -1938
rect 5612 -2040 5646 -2006
rect 5612 -2108 5646 -2074
rect 5612 -2176 5646 -2142
rect 5612 -2244 5646 -2210
rect 5612 -2312 5646 -2278
rect 5612 -2380 5646 -2346
rect 5612 -2448 5646 -2414
rect 5612 -2516 5646 -2482
rect 5612 -2584 5646 -2550
rect 6210 -1874 6244 -1840
rect 6210 -1942 6244 -1908
rect 6210 -2010 6244 -1976
rect 6210 -2078 6244 -2044
rect 6210 -2146 6244 -2112
rect 6210 -2214 6244 -2180
rect 6210 -2282 6244 -2248
rect 6210 -2350 6244 -2316
rect 6210 -2418 6244 -2384
rect 6210 -2486 6244 -2452
rect 6210 -2554 6244 -2520
rect 6808 -1874 6842 -1840
rect 6808 -1942 6842 -1908
rect 6808 -2010 6842 -1976
rect 6808 -2078 6842 -2044
rect 6808 -2146 6842 -2112
rect 6808 -2214 6842 -2180
rect 6808 -2282 6842 -2248
rect 6808 -2350 6842 -2316
rect 6808 -2418 6842 -2384
rect 6808 -2486 6842 -2452
rect 6808 -2554 6842 -2520
rect 7212 -1874 7246 -1840
rect 7212 -1942 7246 -1908
rect 7212 -2010 7246 -1976
rect 7212 -2078 7246 -2044
rect 7212 -2146 7246 -2112
rect 7212 -2214 7246 -2180
rect 7212 -2282 7246 -2248
rect 7212 -2350 7246 -2316
rect 7212 -2418 7246 -2384
rect 7212 -2486 7246 -2452
rect 7212 -2554 7246 -2520
<< locali >>
rect 2478 -1616 2558 -1600
rect 3608 -1824 3642 -1808
rect 3608 -2616 3642 -2600
rect 4012 -1824 4046 -1808
rect 4012 -2616 4046 -2600
rect 4610 -1824 4644 -1808
rect 4610 -2616 4644 -2600
rect 5208 -1824 5242 -1808
rect 5208 -2616 5242 -2600
rect 5612 -1824 5646 -1808
rect 5612 -2616 5646 -2600
rect 6210 -1824 6244 -1808
rect 6210 -2616 6244 -2600
rect 6808 -1824 6842 -1808
rect 6808 -2616 6842 -2600
rect 7212 -1824 7246 -1808
rect 7212 -2616 7246 -2600
rect 2478 -4610 2558 -4494
rect 2672 -3240 2752 -3124
rect 3274 -3240 3354 -3124
rect 3876 -3240 3956 -3124
rect 2672 -6808 2752 -6728
rect 4478 -3240 4558 -3124
rect 3274 -6808 3354 -6728
rect 6034 -3240 6114 -3124
rect 6638 -3240 6718 -3124
rect 5582 -4706 5616 -4690
rect 5582 -5098 5616 -5082
rect 3876 -6808 3956 -6728
rect 4478 -6808 4558 -6728
rect 7242 -3240 7322 -3124
rect 6034 -6808 6114 -6728
rect 7846 -3240 7926 -3124
rect 6638 -6808 6718 -6728
rect 8450 -3240 8530 -3124
rect 7242 -6808 7322 -6728
rect 9054 -3240 9134 -3124
rect 7846 -6808 7926 -6728
rect 8450 -6808 8530 -6728
rect 9054 -6808 9134 -6728
<< viali >>
rect 2478 -1788 2558 -1616
rect 2478 -1888 2558 -1788
rect 2478 -2060 2558 -1888
rect 2478 -2222 2558 -2060
rect 2478 -2394 2558 -2222
rect 2478 -2534 2558 -2394
rect 2478 -2706 2558 -2534
rect 3608 -1840 3642 -1824
rect 3608 -1874 3642 -1840
rect 3608 -1908 3642 -1874
rect 3608 -1942 3642 -1908
rect 3608 -1976 3642 -1942
rect 3608 -2010 3642 -1976
rect 3608 -2044 3642 -2010
rect 3608 -2078 3642 -2044
rect 3608 -2112 3642 -2078
rect 3608 -2146 3642 -2112
rect 3608 -2180 3642 -2146
rect 3608 -2214 3642 -2180
rect 3608 -2248 3642 -2214
rect 3608 -2282 3642 -2248
rect 3608 -2316 3642 -2282
rect 3608 -2350 3642 -2316
rect 3608 -2384 3642 -2350
rect 3608 -2418 3642 -2384
rect 3608 -2452 3642 -2418
rect 3608 -2486 3642 -2452
rect 3608 -2520 3642 -2486
rect 3608 -2554 3642 -2520
rect 3608 -2600 3642 -2554
rect 4012 -1840 4046 -1824
rect 4012 -1874 4046 -1840
rect 4012 -1908 4046 -1874
rect 4012 -1942 4046 -1908
rect 4012 -1976 4046 -1942
rect 4012 -2010 4046 -1976
rect 4012 -2044 4046 -2010
rect 4012 -2078 4046 -2044
rect 4012 -2112 4046 -2078
rect 4012 -2146 4046 -2112
rect 4012 -2180 4046 -2146
rect 4012 -2214 4046 -2180
rect 4012 -2248 4046 -2214
rect 4012 -2282 4046 -2248
rect 4012 -2316 4046 -2282
rect 4012 -2350 4046 -2316
rect 4012 -2384 4046 -2350
rect 4012 -2418 4046 -2384
rect 4012 -2452 4046 -2418
rect 4012 -2486 4046 -2452
rect 4012 -2520 4046 -2486
rect 4012 -2554 4046 -2520
rect 4012 -2600 4046 -2554
rect 4610 -1840 4644 -1824
rect 4610 -1874 4644 -1840
rect 4610 -1908 4644 -1874
rect 4610 -1942 4644 -1908
rect 4610 -1976 4644 -1942
rect 4610 -2010 4644 -1976
rect 4610 -2044 4644 -2010
rect 4610 -2078 4644 -2044
rect 4610 -2112 4644 -2078
rect 4610 -2146 4644 -2112
rect 4610 -2180 4644 -2146
rect 4610 -2214 4644 -2180
rect 4610 -2248 4644 -2214
rect 4610 -2282 4644 -2248
rect 4610 -2316 4644 -2282
rect 4610 -2350 4644 -2316
rect 4610 -2384 4644 -2350
rect 4610 -2418 4644 -2384
rect 4610 -2452 4644 -2418
rect 4610 -2486 4644 -2452
rect 4610 -2520 4644 -2486
rect 4610 -2554 4644 -2520
rect 4610 -2600 4644 -2554
rect 5208 -1870 5242 -1824
rect 5208 -1904 5242 -1870
rect 5208 -1938 5242 -1904
rect 5208 -1972 5242 -1938
rect 5208 -2006 5242 -1972
rect 5208 -2040 5242 -2006
rect 5208 -2074 5242 -2040
rect 5208 -2108 5242 -2074
rect 5208 -2142 5242 -2108
rect 5208 -2176 5242 -2142
rect 5208 -2210 5242 -2176
rect 5208 -2244 5242 -2210
rect 5208 -2278 5242 -2244
rect 5208 -2312 5242 -2278
rect 5208 -2346 5242 -2312
rect 5208 -2380 5242 -2346
rect 5208 -2414 5242 -2380
rect 5208 -2448 5242 -2414
rect 5208 -2482 5242 -2448
rect 5208 -2516 5242 -2482
rect 5208 -2550 5242 -2516
rect 5208 -2584 5242 -2550
rect 5208 -2600 5242 -2584
rect 5612 -1870 5646 -1824
rect 5612 -1904 5646 -1870
rect 5612 -1938 5646 -1904
rect 5612 -1972 5646 -1938
rect 5612 -2006 5646 -1972
rect 5612 -2040 5646 -2006
rect 5612 -2074 5646 -2040
rect 5612 -2108 5646 -2074
rect 5612 -2142 5646 -2108
rect 5612 -2176 5646 -2142
rect 5612 -2210 5646 -2176
rect 5612 -2244 5646 -2210
rect 5612 -2278 5646 -2244
rect 5612 -2312 5646 -2278
rect 5612 -2346 5646 -2312
rect 5612 -2380 5646 -2346
rect 5612 -2414 5646 -2380
rect 5612 -2448 5646 -2414
rect 5612 -2482 5646 -2448
rect 5612 -2516 5646 -2482
rect 5612 -2550 5646 -2516
rect 5612 -2584 5646 -2550
rect 5612 -2600 5646 -2584
rect 6210 -1840 6244 -1824
rect 6210 -1874 6244 -1840
rect 6210 -1908 6244 -1874
rect 6210 -1942 6244 -1908
rect 6210 -1976 6244 -1942
rect 6210 -2010 6244 -1976
rect 6210 -2044 6244 -2010
rect 6210 -2078 6244 -2044
rect 6210 -2112 6244 -2078
rect 6210 -2146 6244 -2112
rect 6210 -2180 6244 -2146
rect 6210 -2214 6244 -2180
rect 6210 -2248 6244 -2214
rect 6210 -2282 6244 -2248
rect 6210 -2316 6244 -2282
rect 6210 -2350 6244 -2316
rect 6210 -2384 6244 -2350
rect 6210 -2418 6244 -2384
rect 6210 -2452 6244 -2418
rect 6210 -2486 6244 -2452
rect 6210 -2520 6244 -2486
rect 6210 -2554 6244 -2520
rect 6210 -2600 6244 -2554
rect 6808 -1840 6842 -1824
rect 6808 -1874 6842 -1840
rect 6808 -1908 6842 -1874
rect 6808 -1942 6842 -1908
rect 6808 -1976 6842 -1942
rect 6808 -2010 6842 -1976
rect 6808 -2044 6842 -2010
rect 6808 -2078 6842 -2044
rect 6808 -2112 6842 -2078
rect 6808 -2146 6842 -2112
rect 6808 -2180 6842 -2146
rect 6808 -2214 6842 -2180
rect 6808 -2248 6842 -2214
rect 6808 -2282 6842 -2248
rect 6808 -2316 6842 -2282
rect 6808 -2350 6842 -2316
rect 6808 -2384 6842 -2350
rect 6808 -2418 6842 -2384
rect 6808 -2452 6842 -2418
rect 6808 -2486 6842 -2452
rect 6808 -2520 6842 -2486
rect 6808 -2554 6842 -2520
rect 6808 -2600 6842 -2554
rect 7212 -1840 7246 -1824
rect 7212 -1874 7246 -1840
rect 7212 -1908 7246 -1874
rect 7212 -1942 7246 -1908
rect 7212 -1976 7246 -1942
rect 7212 -2010 7246 -1976
rect 7212 -2044 7246 -2010
rect 7212 -2078 7246 -2044
rect 7212 -2112 7246 -2078
rect 7212 -2146 7246 -2112
rect 7212 -2180 7246 -2146
rect 7212 -2214 7246 -2180
rect 7212 -2248 7246 -2214
rect 7212 -2282 7246 -2248
rect 7212 -2316 7246 -2282
rect 7212 -2350 7246 -2316
rect 7212 -2384 7246 -2350
rect 7212 -2418 7246 -2384
rect 7212 -2452 7246 -2418
rect 7212 -2486 7246 -2452
rect 7212 -2520 7246 -2486
rect 7212 -2554 7246 -2520
rect 7212 -2600 7246 -2554
rect 2478 -2840 2558 -2706
rect 2478 -3012 2558 -2840
rect 2478 -3098 2558 -3012
rect 2478 -3270 2558 -3098
rect 2478 -3370 2558 -3270
rect 2478 -3542 2558 -3370
rect 2478 -3704 2558 -3542
rect 2478 -3876 2558 -3704
rect 2478 -4016 2558 -3876
rect 2478 -4188 2558 -4016
rect 2478 -4322 2558 -4188
rect 2478 -4494 2558 -4322
rect 2672 -3412 2752 -3240
rect 2672 -3512 2752 -3412
rect 2672 -3684 2752 -3512
rect 2672 -3822 2752 -3684
rect 2672 -3994 2752 -3822
rect 2672 -4094 2752 -3994
rect 2672 -4266 2752 -4094
rect 2672 -4428 2752 -4266
rect 2672 -4600 2752 -4428
rect 2672 -4740 2752 -4600
rect 2672 -4912 2752 -4740
rect 2672 -5046 2752 -4912
rect 2672 -5218 2752 -5046
rect 2672 -5332 2752 -5218
rect 2672 -5504 2752 -5332
rect 2672 -5604 2752 -5504
rect 2672 -5776 2752 -5604
rect 2672 -5938 2752 -5776
rect 2672 -6110 2752 -5938
rect 2672 -6250 2752 -6110
rect 2672 -6422 2752 -6250
rect 3274 -3412 3354 -3240
rect 3274 -3512 3354 -3412
rect 3274 -3684 3354 -3512
rect 3486 -3544 3744 -3136
rect 3876 -3412 3956 -3240
rect 3876 -3512 3956 -3412
rect 3274 -3822 3354 -3684
rect 3274 -3994 3354 -3822
rect 3274 -4094 3354 -3994
rect 3274 -4266 3354 -4094
rect 3274 -4428 3354 -4266
rect 3274 -4600 3354 -4428
rect 3274 -4740 3354 -4600
rect 3274 -4912 3354 -4740
rect 3274 -5046 3354 -4912
rect 3274 -5218 3354 -5046
rect 3274 -5332 3354 -5218
rect 3274 -5504 3354 -5332
rect 3274 -5604 3354 -5504
rect 3274 -5776 3354 -5604
rect 3274 -5938 3354 -5776
rect 3274 -6110 3354 -5938
rect 3274 -6250 3354 -6110
rect 2672 -6556 2752 -6422
rect 2672 -6728 2752 -6556
rect 2884 -6796 3142 -6388
rect 3274 -6422 3354 -6250
rect 3876 -3684 3956 -3512
rect 4088 -3544 4346 -3136
rect 4478 -3412 4558 -3240
rect 4478 -3512 4558 -3412
rect 3876 -3822 3956 -3684
rect 3876 -3994 3956 -3822
rect 3876 -4094 3956 -3994
rect 3876 -4266 3956 -4094
rect 3876 -4428 3956 -4266
rect 3876 -4600 3956 -4428
rect 3876 -4740 3956 -4600
rect 3876 -4912 3956 -4740
rect 3876 -5046 3956 -4912
rect 3876 -5218 3956 -5046
rect 3876 -5332 3956 -5218
rect 3876 -5504 3956 -5332
rect 3876 -5604 3956 -5504
rect 3876 -5776 3956 -5604
rect 3876 -5938 3956 -5776
rect 3876 -6110 3956 -5938
rect 3876 -6250 3956 -6110
rect 3274 -6556 3354 -6422
rect 3274 -6728 3354 -6556
rect 3486 -6796 3744 -6388
rect 3876 -6422 3956 -6250
rect 4478 -3684 4558 -3512
rect 4692 -3544 4950 -3136
rect 6034 -3412 6114 -3240
rect 6034 -3512 6114 -3412
rect 4478 -3822 4558 -3684
rect 4478 -3994 4558 -3822
rect 4478 -4094 4558 -3994
rect 4478 -4266 4558 -4094
rect 4478 -4428 4558 -4266
rect 4478 -4600 4558 -4428
rect 4478 -4740 4558 -4600
rect 6034 -3684 6114 -3512
rect 6248 -3544 6506 -3136
rect 6638 -3412 6718 -3240
rect 6638 -3512 6718 -3412
rect 6034 -3822 6114 -3684
rect 6034 -3994 6114 -3822
rect 6034 -4094 6114 -3994
rect 6034 -4266 6114 -4094
rect 6034 -4428 6114 -4266
rect 6034 -4600 6114 -4428
rect 4478 -4912 4558 -4740
rect 4478 -5046 4558 -4912
rect 4478 -5218 4558 -5046
rect 5582 -4760 5616 -4706
rect 5582 -4794 5616 -4760
rect 5582 -4828 5616 -4794
rect 5582 -4862 5616 -4828
rect 5582 -4896 5616 -4862
rect 5582 -4930 5616 -4896
rect 5582 -4964 5616 -4930
rect 5582 -4998 5616 -4964
rect 5582 -5032 5616 -4998
rect 5582 -5066 5616 -5032
rect 5582 -5082 5616 -5066
rect 6034 -4740 6114 -4600
rect 6034 -4912 6114 -4740
rect 6034 -5046 6114 -4912
rect 4478 -5332 4558 -5218
rect 4478 -5504 4558 -5332
rect 4478 -5604 4558 -5504
rect 4478 -5776 4558 -5604
rect 4478 -5938 4558 -5776
rect 4478 -6110 4558 -5938
rect 4478 -6250 4558 -6110
rect 3876 -6556 3956 -6422
rect 3876 -6728 3956 -6556
rect 4088 -6796 4346 -6388
rect 4478 -6422 4558 -6250
rect 6034 -5218 6114 -5046
rect 6034 -5332 6114 -5218
rect 6034 -5504 6114 -5332
rect 6034 -5604 6114 -5504
rect 6034 -5776 6114 -5604
rect 6034 -5938 6114 -5776
rect 6034 -6110 6114 -5938
rect 6034 -6250 6114 -6110
rect 4478 -6556 4558 -6422
rect 4478 -6728 4558 -6556
rect 4692 -6796 4950 -6388
rect 6034 -6422 6114 -6250
rect 6638 -3684 6718 -3512
rect 6852 -3544 7110 -3136
rect 7242 -3412 7322 -3240
rect 7242 -3512 7322 -3412
rect 6638 -3822 6718 -3684
rect 6638 -3994 6718 -3822
rect 6638 -4094 6718 -3994
rect 6638 -4266 6718 -4094
rect 6638 -4428 6718 -4266
rect 6638 -4600 6718 -4428
rect 6638 -4740 6718 -4600
rect 6638 -4912 6718 -4740
rect 6638 -5046 6718 -4912
rect 6638 -5218 6718 -5046
rect 6638 -5332 6718 -5218
rect 6638 -5504 6718 -5332
rect 6638 -5604 6718 -5504
rect 6638 -5776 6718 -5604
rect 6638 -5938 6718 -5776
rect 6638 -6110 6718 -5938
rect 6638 -6250 6718 -6110
rect 6034 -6556 6114 -6422
rect 6034 -6728 6114 -6556
rect 6248 -6796 6506 -6388
rect 6638 -6422 6718 -6250
rect 7242 -3684 7322 -3512
rect 7456 -3544 7714 -3136
rect 7846 -3412 7926 -3240
rect 7846 -3512 7926 -3412
rect 7242 -3822 7322 -3684
rect 7242 -3994 7322 -3822
rect 7242 -4094 7322 -3994
rect 7242 -4266 7322 -4094
rect 7242 -4428 7322 -4266
rect 7242 -4600 7322 -4428
rect 7242 -4740 7322 -4600
rect 7242 -4912 7322 -4740
rect 7242 -5046 7322 -4912
rect 7242 -5218 7322 -5046
rect 7242 -5332 7322 -5218
rect 7242 -5504 7322 -5332
rect 7242 -5604 7322 -5504
rect 7242 -5776 7322 -5604
rect 7242 -5938 7322 -5776
rect 7242 -6110 7322 -5938
rect 7242 -6250 7322 -6110
rect 6638 -6556 6718 -6422
rect 6638 -6728 6718 -6556
rect 6852 -6796 7110 -6388
rect 7242 -6422 7322 -6250
rect 7846 -3684 7926 -3512
rect 8060 -3544 8318 -3136
rect 8450 -3412 8530 -3240
rect 8450 -3512 8530 -3412
rect 7846 -3822 7926 -3684
rect 7846 -3994 7926 -3822
rect 7846 -4094 7926 -3994
rect 7846 -4266 7926 -4094
rect 7846 -4428 7926 -4266
rect 7846 -4600 7926 -4428
rect 7846 -4740 7926 -4600
rect 7846 -4912 7926 -4740
rect 7846 -5046 7926 -4912
rect 7846 -5218 7926 -5046
rect 7846 -5332 7926 -5218
rect 7846 -5504 7926 -5332
rect 7846 -5604 7926 -5504
rect 7846 -5776 7926 -5604
rect 7846 -5938 7926 -5776
rect 7846 -6110 7926 -5938
rect 7846 -6250 7926 -6110
rect 7242 -6556 7322 -6422
rect 7242 -6728 7322 -6556
rect 7456 -6796 7714 -6388
rect 7846 -6422 7926 -6250
rect 8450 -3684 8530 -3512
rect 8664 -3544 8922 -3136
rect 9054 -3412 9134 -3240
rect 9054 -3512 9134 -3412
rect 8450 -3822 8530 -3684
rect 8450 -3994 8530 -3822
rect 8450 -4094 8530 -3994
rect 8450 -4266 8530 -4094
rect 8450 -4428 8530 -4266
rect 8450 -4600 8530 -4428
rect 8450 -4740 8530 -4600
rect 8450 -4912 8530 -4740
rect 8450 -5046 8530 -4912
rect 8450 -5218 8530 -5046
rect 8450 -5332 8530 -5218
rect 8450 -5504 8530 -5332
rect 8450 -5604 8530 -5504
rect 8450 -5776 8530 -5604
rect 8450 -5938 8530 -5776
rect 8450 -6110 8530 -5938
rect 8450 -6250 8530 -6110
rect 7846 -6556 7926 -6422
rect 7846 -6728 7926 -6556
rect 8060 -6796 8318 -6388
rect 8450 -6422 8530 -6250
rect 9054 -3684 9134 -3512
rect 9054 -3822 9134 -3684
rect 9054 -3994 9134 -3822
rect 9054 -4094 9134 -3994
rect 9054 -4266 9134 -4094
rect 9054 -4428 9134 -4266
rect 9054 -4600 9134 -4428
rect 9054 -4740 9134 -4600
rect 9054 -4912 9134 -4740
rect 9054 -5046 9134 -4912
rect 9054 -5218 9134 -5046
rect 9054 -5332 9134 -5218
rect 9054 -5504 9134 -5332
rect 9054 -5604 9134 -5504
rect 9054 -5776 9134 -5604
rect 9054 -5938 9134 -5776
rect 9054 -6110 9134 -5938
rect 9054 -6250 9134 -6110
rect 8450 -6556 8530 -6422
rect 8450 -6728 8530 -6556
rect 8664 -6796 8922 -6388
rect 9054 -6422 9134 -6250
rect 9054 -6556 9134 -6422
rect 9054 -6728 9134 -6556
rect 9268 -6796 9526 -6388
<< metal1 >>
rect 1216 -904 2354 -898
rect 1216 -1836 2354 -1354
rect 3592 -904 3704 -898
rect 1212 -3770 2354 -1836
rect 2472 -1616 2564 -1600
rect 2472 -4494 2478 -1616
rect 2558 -2430 2564 -1616
rect 3592 -1812 3704 -1354
rect 3996 -904 4108 -898
rect 3732 -1688 3738 -1576
rect 3962 -1688 3968 -1576
rect 3732 -1694 3968 -1688
rect 3732 -1772 3794 -1694
rect 3860 -1772 3922 -1694
rect 3996 -1812 4108 -1354
rect 4592 -904 4650 -898
rect 4136 -1778 4316 -1688
rect 3592 -1824 3722 -1812
rect 2558 -3124 2582 -2430
rect 3592 -2600 3608 -1824
rect 3642 -2600 3722 -1824
rect 3592 -2612 3722 -2600
rect 3800 -1824 3852 -1818
rect 3800 -2606 3852 -2600
rect 3932 -1824 4126 -1812
rect 3932 -2600 4012 -1824
rect 4046 -2600 4126 -1824
rect 3932 -2612 4126 -2600
rect 4208 -2820 4316 -1778
rect 4592 -1824 4650 -1354
rect 5190 -904 5248 -898
rect 4754 -1782 4884 -1724
rect 4592 -2600 4610 -1824
rect 4644 -2600 4650 -1824
rect 4592 -2612 4650 -2600
rect 4678 -2820 4776 -1812
rect 4826 -2674 4884 -1782
rect 5190 -1824 5248 -1354
rect 5606 -904 5664 -898
rect 5332 -1772 5522 -1724
rect 5190 -2600 5208 -1824
rect 5242 -2600 5248 -1824
rect 5190 -2612 5248 -2600
rect 5276 -2674 5334 -1812
rect 4826 -2680 4950 -2674
rect 4826 -2792 4832 -2680
rect 4944 -2792 4950 -2680
rect 4826 -2798 4950 -2792
rect 5210 -2680 5334 -2674
rect 5210 -2792 5216 -2680
rect 5328 -2792 5334 -2680
rect 5210 -2798 5334 -2792
rect 4208 -2826 4332 -2820
rect 4208 -2938 4214 -2826
rect 4326 -2938 4332 -2826
rect 4208 -2944 4332 -2938
rect 4666 -2826 4790 -2820
rect 4666 -2938 4672 -2826
rect 4784 -2938 4790 -2826
rect 4666 -2944 4790 -2938
rect 2558 -3240 2758 -3124
rect 2558 -4494 2672 -3240
rect 2472 -4610 2672 -4494
rect 2480 -6728 2672 -4610
rect 2752 -6728 2758 -3240
rect 2882 -3132 3144 -3124
rect 2882 -3540 2892 -3132
rect 3130 -3540 3144 -3132
rect 3474 -3136 3756 -3124
rect 2882 -3550 3144 -3540
rect 3268 -3240 3360 -3226
rect 2480 -7120 2758 -6728
rect 2872 -6388 3154 -6376
rect 2872 -6796 2884 -6388
rect 3142 -6796 3154 -6388
rect 2872 -6808 3154 -6796
rect 3268 -6728 3274 -3240
rect 3354 -6728 3360 -3240
rect 3474 -3544 3486 -3136
rect 3744 -3544 3756 -3136
rect 3474 -3556 3756 -3544
rect 3870 -3240 3962 -3124
rect 2480 -7576 2758 -7570
rect 2882 -7120 3144 -6808
rect 2882 -7576 3144 -7570
rect 3268 -7120 3360 -6728
rect 3474 -6388 3756 -6376
rect 3474 -6796 3486 -6388
rect 3744 -6796 3756 -6388
rect 3474 -6808 3756 -6796
rect 3870 -6728 3876 -3240
rect 3956 -6728 3962 -3240
rect 4076 -3136 4358 -3124
rect 4076 -3544 4088 -3136
rect 4346 -3544 4358 -3136
rect 4076 -3556 4358 -3544
rect 4472 -3240 4564 -3124
rect 3268 -7576 3360 -7570
rect 3870 -7120 3962 -6728
rect 4076 -6388 4358 -6376
rect 4076 -6796 4088 -6388
rect 4346 -6796 4358 -6388
rect 4076 -6808 4358 -6796
rect 4472 -6728 4478 -3240
rect 4558 -6728 4564 -3240
rect 4680 -3136 4962 -3124
rect 4680 -3544 4692 -3136
rect 4950 -3544 4962 -3136
rect 4680 -3556 4962 -3544
rect 5268 -3298 5332 -3292
rect 5268 -3398 5274 -3298
rect 5326 -3398 5332 -3298
rect 5268 -4694 5332 -3398
rect 5372 -4640 5480 -1772
rect 5520 -2674 5578 -1812
rect 5606 -1824 5664 -1354
rect 6204 -904 6262 -898
rect 5606 -2600 5612 -1824
rect 5646 -2600 5664 -1824
rect 5606 -2612 5664 -2600
rect 5970 -1776 6100 -1718
rect 5970 -2674 6028 -1776
rect 5520 -2680 5644 -2674
rect 5520 -2792 5526 -2680
rect 5638 -2792 5644 -2680
rect 5520 -2798 5644 -2792
rect 5904 -2680 6028 -2674
rect 5904 -2792 5910 -2680
rect 6022 -2792 6028 -2680
rect 5904 -2798 6028 -2792
rect 6098 -2820 6176 -1812
rect 6204 -1824 6262 -1354
rect 6746 -904 6858 -898
rect 6204 -2600 6210 -1824
rect 6244 -2600 6262 -1824
rect 6204 -2612 6262 -2600
rect 6292 -1584 6494 -1576
rect 6292 -1680 6300 -1584
rect 6486 -1680 6494 -1584
rect 6078 -2826 6202 -2820
rect 6078 -2938 6084 -2826
rect 6196 -2938 6202 -2826
rect 6078 -2944 6202 -2938
rect 6292 -3056 6494 -1680
rect 6552 -1780 6718 -1722
rect 6552 -2820 6646 -1780
rect 6746 -1812 6858 -1354
rect 7150 -904 7262 -898
rect 6886 -1576 7122 -1570
rect 6886 -1688 6892 -1576
rect 7116 -1688 7122 -1576
rect 6886 -1694 7122 -1688
rect 6932 -1772 6994 -1694
rect 7060 -1772 7122 -1694
rect 7150 -1812 7262 -1354
rect 6728 -1824 6922 -1812
rect 6728 -2600 6808 -1824
rect 6842 -2600 6922 -1824
rect 6728 -2612 6922 -2600
rect 7000 -1824 7052 -1818
rect 7000 -2606 7052 -2600
rect 7132 -1824 7262 -1812
rect 7132 -2600 7212 -1824
rect 7246 -2600 7262 -1824
rect 7132 -2612 7262 -2600
rect 9266 -904 9528 -898
rect 6932 -2710 7122 -2652
rect 6522 -2826 6646 -2820
rect 6522 -2938 6528 -2826
rect 6640 -2938 6646 -2826
rect 6522 -2944 6646 -2938
rect 6028 -3240 6120 -3124
rect 5394 -4644 5452 -4640
rect 5268 -5094 5350 -4694
rect 5502 -4704 5622 -4694
rect 5502 -5084 5516 -4704
rect 5610 -4706 5622 -4704
rect 5616 -5082 5622 -4706
rect 5610 -5084 5622 -5082
rect 5502 -5094 5622 -5084
rect 3870 -7576 3962 -7570
rect 4472 -7120 4564 -6728
rect 4680 -6388 4962 -6376
rect 4680 -6796 4692 -6388
rect 4950 -6796 4962 -6388
rect 4680 -6808 4962 -6796
rect 5372 -6388 5480 -5172
rect 5372 -6796 5378 -6388
rect 5474 -6796 5480 -6388
rect 5372 -6802 5480 -6796
rect 6028 -6728 6034 -3240
rect 6114 -6728 6120 -3240
rect 6236 -3136 6518 -3056
rect 6236 -3544 6248 -3136
rect 6506 -3544 6518 -3136
rect 6236 -3556 6518 -3544
rect 6632 -3240 6724 -3124
rect 4472 -7576 4564 -7570
rect 6028 -7120 6120 -6728
rect 6236 -6388 6518 -6376
rect 6236 -6796 6248 -6388
rect 6506 -6796 6518 -6388
rect 6236 -6808 6518 -6796
rect 6632 -6728 6638 -3240
rect 6718 -6728 6724 -3240
rect 6840 -3136 7122 -3124
rect 6840 -3544 6852 -3136
rect 7110 -3544 7122 -3136
rect 6840 -3556 7122 -3544
rect 7236 -3240 7328 -3124
rect 6028 -7576 6120 -7570
rect 6632 -7120 6724 -6728
rect 6840 -6388 7122 -6376
rect 6840 -6796 6852 -6388
rect 7110 -6796 7122 -6388
rect 6840 -6808 7122 -6796
rect 7236 -6728 7242 -3240
rect 7322 -6728 7328 -3240
rect 7444 -3136 7726 -3124
rect 7444 -3544 7456 -3136
rect 7714 -3544 7726 -3136
rect 7444 -3556 7726 -3544
rect 7840 -3240 7932 -3124
rect 6632 -7576 6724 -7570
rect 7236 -7120 7328 -6728
rect 7444 -6388 7726 -6376
rect 7444 -6796 7456 -6388
rect 7714 -6796 7726 -6388
rect 7444 -6808 7726 -6796
rect 7840 -6728 7846 -3240
rect 7926 -6728 7932 -3240
rect 8048 -3136 8330 -3124
rect 8048 -3544 8060 -3136
rect 8318 -3544 8330 -3136
rect 8048 -3556 8330 -3544
rect 8444 -3240 8536 -3124
rect 7236 -7576 7328 -7570
rect 7840 -7120 7932 -6728
rect 8048 -6388 8330 -6376
rect 8048 -6796 8060 -6388
rect 8318 -6796 8330 -6388
rect 8048 -6808 8330 -6796
rect 8444 -6728 8450 -3240
rect 8530 -6728 8536 -3240
rect 8652 -3136 8934 -3124
rect 8652 -3544 8664 -3136
rect 8922 -3544 8934 -3136
rect 8652 -3556 8934 -3544
rect 9048 -3240 9140 -3124
rect 7840 -7576 7932 -7570
rect 8444 -7120 8536 -6728
rect 8652 -6388 8934 -6376
rect 8652 -6796 8664 -6388
rect 8922 -6796 8934 -6388
rect 8652 -6808 8934 -6796
rect 9048 -6728 9054 -3240
rect 9134 -6728 9140 -3240
rect 9266 -3550 9528 -1354
rect 8444 -7576 8536 -7570
rect 9048 -7120 9140 -6728
rect 9256 -6388 9538 -6376
rect 9256 -6796 9268 -6388
rect 9526 -6796 9538 -6388
rect 9256 -6808 9538 -6796
rect 9048 -7576 9140 -7570
<< via1 >>
rect 1216 -1354 2354 -904
rect 3592 -1354 3704 -904
rect 1228 -4592 2342 -4196
rect 3996 -1354 4108 -904
rect 3738 -1688 3962 -1576
rect 4592 -1354 4650 -904
rect 3800 -2600 3852 -1824
rect 5190 -1354 5248 -904
rect 5606 -1354 5664 -904
rect 4832 -2792 4944 -2680
rect 5216 -2792 5328 -2680
rect 4214 -2938 4326 -2826
rect 4672 -2938 4784 -2826
rect 2892 -3540 3130 -3132
rect 2884 -6796 3142 -6388
rect 3486 -3544 3744 -3136
rect 2480 -7570 2758 -7120
rect 2882 -7570 3144 -7120
rect 3486 -6796 3744 -6388
rect 3890 -4804 3942 -4028
rect 3890 -5592 3942 -4816
rect 4088 -3544 4346 -3136
rect 3268 -7570 3360 -7120
rect 4088 -6796 4346 -6388
rect 4692 -3544 4950 -3136
rect 5274 -3398 5326 -3298
rect 6204 -1354 6262 -904
rect 5526 -2792 5638 -2680
rect 5910 -2792 6022 -2680
rect 6746 -1354 6858 -904
rect 6300 -1680 6486 -1584
rect 6084 -2938 6196 -2826
rect 7150 -1354 7262 -904
rect 6892 -1688 7116 -1576
rect 7000 -2600 7052 -1824
rect 9266 -1354 9528 -904
rect 6528 -2938 6640 -2826
rect 5516 -4706 5610 -4704
rect 5516 -5082 5582 -4706
rect 5582 -5082 5610 -4706
rect 5516 -5084 5610 -5082
rect 3870 -7570 3962 -7120
rect 4692 -6796 4950 -6388
rect 5378 -6796 5474 -6388
rect 6038 -5088 6110 -4702
rect 6248 -3544 6506 -3136
rect 4472 -7570 4564 -7120
rect 6248 -6796 6506 -6388
rect 6852 -3544 7110 -3136
rect 6028 -7570 6120 -7120
rect 6852 -6796 7110 -6388
rect 7256 -4804 7308 -4028
rect 7256 -5592 7308 -4816
rect 7456 -3544 7714 -3136
rect 6632 -7570 6724 -7120
rect 7456 -6796 7714 -6388
rect 8060 -3544 8318 -3136
rect 7236 -7570 7328 -7120
rect 8060 -6796 8318 -6388
rect 8664 -3544 8922 -3136
rect 7840 -7570 7932 -7120
rect 8664 -6796 8922 -6388
rect 8444 -7570 8536 -7120
rect 9268 -6796 9526 -6388
rect 9048 -7570 9140 -7120
<< metal2 >>
rect 658 -904 9804 -892
rect 658 -1354 1216 -904
rect 2354 -1354 3592 -904
rect 3704 -1354 3996 -904
rect 4108 -1354 4592 -904
rect 4650 -1354 5190 -904
rect 5248 -1354 5606 -904
rect 5664 -1354 6204 -904
rect 6262 -1354 6746 -904
rect 6858 -1354 7150 -904
rect 7262 -1354 9266 -904
rect 9528 -1354 9804 -904
rect 658 -1360 9804 -1354
rect 6886 -1576 7122 -1570
rect 3732 -1688 3738 -1576
rect 3962 -1584 6892 -1576
rect 3962 -1680 6300 -1584
rect 6486 -1680 6892 -1584
rect 3962 -1688 6892 -1680
rect 7116 -1688 7122 -1576
rect 3732 -1694 3968 -1688
rect 6886 -1694 7122 -1688
rect 3798 -1824 3854 -1814
rect 3798 -2610 3854 -2600
rect 6998 -1824 7054 -1814
rect 6998 -2610 7054 -2600
rect 4826 -2680 4950 -2674
rect 5210 -2680 5334 -2674
rect 5520 -2680 5644 -2674
rect 5904 -2680 6028 -2674
rect 4826 -2792 4832 -2680
rect 4944 -2792 5216 -2680
rect 5328 -2792 5526 -2680
rect 5638 -2792 5910 -2680
rect 6022 -2792 6028 -2680
rect 4826 -2798 4950 -2792
rect 5210 -2798 5334 -2792
rect 5520 -2798 5644 -2792
rect 5904 -2798 6028 -2792
rect 4208 -2826 4332 -2820
rect 4666 -2826 4790 -2820
rect 6078 -2826 6202 -2820
rect 6522 -2826 6646 -2820
rect 4208 -2938 4214 -2826
rect 4326 -2938 4672 -2826
rect 4784 -2938 6084 -2826
rect 6196 -2938 6528 -2826
rect 6640 -2938 6646 -2826
rect 4208 -2944 4332 -2938
rect 4666 -2944 4790 -2938
rect 6078 -2944 6202 -2938
rect 6522 -2944 6646 -2938
rect 2884 -3132 3750 -3130
rect 2884 -3540 2892 -3132
rect 3130 -3136 3750 -3132
rect 3130 -3540 3486 -3136
rect 2884 -3544 3486 -3540
rect 3744 -3544 3750 -3136
rect 2884 -3550 3750 -3544
rect 4082 -3136 4956 -3130
rect 4082 -3544 4088 -3136
rect 4346 -3544 4692 -3136
rect 4950 -3544 4956 -3136
rect 6242 -3136 6512 -3130
rect 6242 -3292 6248 -3136
rect 5268 -3298 6248 -3292
rect 5268 -3398 5274 -3298
rect 5326 -3398 6248 -3298
rect 5268 -3404 6248 -3398
rect 4082 -3550 4956 -3544
rect 6242 -3544 6248 -3404
rect 6506 -3544 6512 -3136
rect 6242 -3550 6512 -3544
rect 6846 -3136 7720 -3130
rect 6846 -3544 6852 -3136
rect 7110 -3544 7456 -3136
rect 7714 -3544 7720 -3136
rect 6846 -3550 7720 -3544
rect 8054 -3136 8928 -3130
rect 8054 -3544 8060 -3136
rect 8318 -3544 8664 -3136
rect 8922 -3544 8928 -3136
rect 8054 -3550 8928 -3544
rect 3888 -4028 3944 -4018
rect 660 -4190 2354 -4180
rect 660 -6966 670 -4190
rect 1186 -4196 2354 -4190
rect 1186 -4592 1228 -4196
rect 2342 -4592 2354 -4196
rect 1186 -4610 2354 -4592
rect 7254 -4028 7310 -4018
rect 5504 -4702 6120 -4694
rect 5504 -4704 6038 -4702
rect 5504 -5084 5516 -4704
rect 5610 -5084 6038 -4704
rect 5504 -5088 6038 -5084
rect 6110 -5088 6120 -4702
rect 5504 -5092 6120 -5088
rect 3888 -5602 3944 -5592
rect 7254 -5602 7310 -5592
rect 2878 -6388 3156 -6382
rect 2878 -6796 2884 -6388
rect 3142 -6796 3156 -6388
rect 2878 -6802 3156 -6796
rect 3480 -6388 4352 -6382
rect 3480 -6796 3486 -6388
rect 3744 -6796 4088 -6388
rect 4346 -6796 4352 -6388
rect 3480 -6802 4352 -6796
rect 4686 -6388 5480 -6382
rect 4686 -6796 4692 -6388
rect 4950 -6796 5378 -6388
rect 5474 -6796 5480 -6388
rect 4686 -6802 5480 -6796
rect 6242 -6388 7116 -6382
rect 6242 -6796 6248 -6388
rect 6506 -6796 6852 -6388
rect 7110 -6796 7116 -6388
rect 6242 -6802 7116 -6796
rect 7450 -6388 8324 -6382
rect 7450 -6796 7456 -6388
rect 7714 -6796 8060 -6388
rect 8318 -6796 8324 -6388
rect 7450 -6802 8324 -6796
rect 8658 -6388 9532 -6382
rect 8658 -6796 8664 -6388
rect 8922 -6796 9268 -6388
rect 9526 -6796 9532 -6388
rect 8658 -6802 9532 -6796
rect 660 -6976 1186 -6966
rect 658 -7120 9804 -7114
rect 658 -7570 2480 -7120
rect 2758 -7570 2882 -7120
rect 3144 -7570 3268 -7120
rect 3360 -7570 3870 -7120
rect 3962 -7570 4472 -7120
rect 4564 -7570 6028 -7120
rect 6120 -7570 6632 -7120
rect 6724 -7570 7236 -7120
rect 7328 -7570 7840 -7120
rect 7932 -7570 8444 -7120
rect 8536 -7570 9048 -7120
rect 9140 -7570 9804 -7120
rect 658 -7582 9804 -7570
<< via2 >>
rect 3798 -2600 3800 -1824
rect 3800 -2600 3852 -1824
rect 3852 -2600 3854 -1824
rect 6998 -2600 7000 -1824
rect 7000 -2600 7052 -1824
rect 7052 -2600 7054 -1824
rect 670 -6966 1186 -4190
rect 1228 -4592 2342 -4196
rect 3888 -4804 3890 -4028
rect 3890 -4804 3942 -4028
rect 3942 -4804 3944 -4028
rect 3888 -4816 3944 -4804
rect 3888 -5592 3890 -4816
rect 3890 -5592 3942 -4816
rect 3942 -5592 3944 -4816
rect 7254 -4804 7256 -4028
rect 7256 -4804 7308 -4028
rect 7308 -4804 7310 -4028
rect 7254 -4816 7310 -4804
rect 7254 -5592 7256 -4816
rect 7256 -5592 7308 -4816
rect 7308 -5592 7310 -4816
<< metal3 >>
rect 3792 -1824 3860 -1818
rect 3792 -2600 3798 -1824
rect 3854 -2600 3860 -1824
rect 3792 -2886 3860 -2600
rect 6992 -1824 7060 -1818
rect 6992 -2600 6998 -1824
rect 7054 -2600 7060 -1824
rect 6992 -2732 7060 -2600
rect 6992 -2800 7316 -2732
rect 3792 -2954 3950 -2886
rect 3882 -4028 3950 -2954
rect 658 -4190 1198 -4178
rect 658 -6966 670 -4190
rect 1186 -4196 2348 -4190
rect 1186 -4592 1228 -4196
rect 2342 -4592 2348 -4196
rect 1186 -6966 2348 -4592
rect 3882 -5592 3888 -4028
rect 3944 -5592 3950 -4028
rect 3882 -5598 3950 -5592
rect 7248 -4028 7316 -2800
rect 7248 -5592 7254 -4028
rect 7310 -5592 7316 -4028
rect 7248 -5598 7316 -5592
rect 658 -6978 2348 -6966
use sky130_fd_pr__nfet_01v8_lvt_BNLWPS  M4
timestamp 1680390383
transform 1 0 5426 0 1 -4894
box -128 -288 128 288
use sky130_fd_pr__pfet_01v8_lvt_73XLH3  M11
timestamp 1680972802
transform -1 0 4167 0 -1 -2176
box -129 -464 129 498
use sky130_fd_pr__pfet_01v8_lvt_73XLH3  M12
timestamp 1680972802
transform 1 0 6687 0 -1 -2176
box -129 -464 129 498
use sky130_fd_pr__pfet_01v8_lvt_73XLH3  M21
timestamp 1680972802
transform -1 0 4785 0 -1 -2176
box -129 -464 129 498
use sky130_fd_pr__pfet_01v8_lvt_73XLH3  M22
timestamp 1680972802
transform 1 0 6069 0 -1 -2176
box -129 -464 129 498
use sky130_fd_pr__pfet_01v8_lvt_M2XLH9  M31
timestamp 1680985943
transform 1 0 5363 0 1 -2176
box -129 -498 129 464
use sky130_fd_pr__pfet_01v8_lvt_M2XLH9  M32
timestamp 1680985943
transform -1 0 5491 0 1 -2176
box -129 -498 129 464
use sky130_fd_pr__pfet_01v8_lvt_73XLH3  M51
timestamp 1680972802
transform -1 0 3763 0 -1 -2176
box -129 -464 129 498
use sky130_fd_pr__pfet_01v8_lvt_73XLH3  M52
timestamp 1680972802
transform 1 0 3891 0 -1 -2176
box -129 -464 129 498
use sky130_fd_pr__pfet_01v8_lvt_4QXLH3  M53
timestamp 1680390383
transform -1 0 6963 0 -1 -2212
box -129 -500 129 500
use sky130_fd_pr__pfet_01v8_lvt_4QXLH3  M54
timestamp 1680390383
transform 1 0 7091 0 -1 -2212
box -129 -500 129 500
use sky130_fd_pr__res_xhigh_po_5p73_J6N8L2  XR2
timestamp 1681965435
transform -1 0 1785 0 1 -4128
box -575 -482 575 482
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR21
timestamp 1680448829
transform 1 0 3013 0 -1 -4966
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR22
timestamp 1680448829
transform 1 0 3615 0 1 -4966
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR23
timestamp 1680448829
transform 1 0 4217 0 -1 -4966
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR24
timestamp 1680448829
transform 1 0 4821 0 1 -4966
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR31
timestamp 1680448829
transform 1 0 6377 0 1 -4966
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR32
timestamp 1680448829
transform 1 0 6981 0 -1 -4966
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR33
timestamp 1680448829
transform 1 0 7585 0 1 -4966
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR34
timestamp 1680448829
transform 1 0 8189 0 -1 -4966
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR35
timestamp 1680448829
transform 1 0 8793 0 1 -4966
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR36
timestamp 1680448829
transform 1 0 9397 0 -1 -4966
box -143 -1842 143 1842
<< labels >>
flabel metal3 658 -6978 1198 -4178 0 FreeMono 1280 90 0 0 vrec
port 0 nsew
flabel metal2 658 -1360 9804 -892 0 FreeMono 1280 0 0 0 vdd
port 1 nsew
flabel metal2 658 -7582 9804 -7114 0 FreeMono 2400 0 0 0 vss
port 2 nsew
<< end >>
