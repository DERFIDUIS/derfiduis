magic
tech sky130A
magscale 1 2
timestamp 1681683204
<< error_p >>
rect -29 -311 29 -305
rect -29 -345 -17 -311
rect -29 -351 29 -345
<< nwell >>
rect -112 -364 112 398
<< pmos >>
rect -18 -264 18 336
<< pdiff >>
rect -76 324 -18 336
rect -76 -252 -64 324
rect -30 -252 -18 324
rect -76 -264 -18 -252
rect 18 324 76 336
rect 18 -252 30 324
rect 64 -252 76 324
rect 18 -264 76 -252
<< pdiffc >>
rect -64 -252 -30 324
rect 30 -252 64 324
<< poly >>
rect -18 336 18 362
rect -18 -295 18 -264
rect -33 -311 33 -295
rect -33 -345 -17 -311
rect 17 -345 33 -311
rect -33 -361 33 -345
<< polycont >>
rect -17 -345 17 -311
<< locali >>
rect -64 324 -30 340
rect -64 -268 -30 -252
rect 30 324 64 340
rect 30 -268 64 -252
rect -33 -345 -17 -311
rect 17 -345 33 -311
<< viali >>
rect -64 -252 -30 324
rect 30 -252 64 324
rect -17 -345 17 -311
<< metal1 >>
rect -70 324 -24 336
rect -70 -252 -64 324
rect -30 -252 -24 324
rect -70 -264 -24 -252
rect 24 324 70 336
rect 24 -252 30 324
rect 64 -252 70 324
rect 24 -264 70 -252
rect -29 -311 29 -305
rect -29 -345 -17 -311
rect 17 -345 29 -311
rect -29 -351 29 -345
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.0 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
