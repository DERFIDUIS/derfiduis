magic
tech sky130A
timestamp 1681769388
<< metal1 >>
rect 9537 17044 9649 17048
rect 9537 16864 9541 17044
rect 9645 16864 9649 17044
rect 9537 16450 9649 16864
rect 12450 17044 12562 17048
rect 12450 16864 12454 17044
rect 12558 16864 12562 17044
rect 12450 16488 12562 16864
rect 12750 16597 12828 17244
rect 9558 15803 9628 16450
rect 12450 15952 12454 16488
rect 12558 15952 12562 16488
rect 12450 15948 12562 15952
rect 9550 14274 9662 15695
rect 9550 14094 9554 14274
rect 9658 14094 9662 14274
rect 9550 14090 9662 14094
rect 12798 14274 12910 15566
rect 12798 14094 12802 14274
rect 12906 14094 12910 14274
rect 12798 14090 12910 14094
<< via1 >>
rect 9541 16864 9645 17044
rect 12454 16864 12558 17044
rect 12454 15952 12558 16488
rect 9554 14094 9658 14274
rect 12802 14094 12906 14274
<< metal2 >>
rect 9567 17574 9610 17798
rect 12767 17574 12810 17798
rect 9537 17044 12562 17048
rect 9537 16864 9541 17044
rect 9645 16864 12454 17044
rect 12558 16864 12562 17044
rect 9537 16860 12562 16864
rect 12562 16491 12802 16492
rect 12450 16488 12802 16491
rect 12450 15952 12454 16488
rect 12558 15952 12802 16488
rect 12450 15948 12802 15952
rect 9550 14274 12910 14278
rect 9550 14094 9554 14274
rect 9658 14094 12802 14274
rect 12906 14094 12910 14274
rect 9550 14090 12910 14094
rect 9568 13631 9611 13855
rect 12774 13631 13074 13855
use BGR_lvt  BGR_lvt_0
timestamp 1681761095
transform 1 0 3778 0 1 18918
box 573 -5287 5793 -1120
use OPAMP_lvt_PMOS  OPAMP_lvt_PMOS_0
timestamp 1681766136
transform 1 0 7940 0 1 16179
box 1668 -2548 4836 1619
use current_source  current_source_0
timestamp 1681769244
transform 1 0 12795 0 1 17814
box 2 -4183 3419 -16
<< end >>
