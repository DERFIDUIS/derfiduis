magic
tech sky130A
magscale 1 2
timestamp 1681051265
<< error_p >>
rect -29 -507 29 -501
rect -29 -541 -17 -507
rect -29 -547 29 -541
<< nmoslvt >>
rect -18 -469 18 531
<< ndiff >>
rect -76 519 -18 531
rect -76 -457 -64 519
rect -30 -457 -18 519
rect -76 -469 -18 -457
rect 18 519 76 531
rect 18 -457 30 519
rect 64 -457 76 519
rect 18 -469 76 -457
<< ndiffc >>
rect -64 -457 -30 519
rect 30 -457 64 519
<< poly >>
rect -18 531 18 557
rect -18 -491 18 -469
rect -33 -507 33 -491
rect -33 -541 -17 -507
rect 17 -541 33 -507
rect -33 -557 33 -541
<< polycont >>
rect -17 -541 17 -507
<< locali >>
rect -64 519 -30 535
rect -64 -473 -30 -457
rect 30 519 64 535
rect 30 -473 64 -457
rect -33 -541 -17 -507
rect 17 -541 33 -507
<< viali >>
rect -64 -457 -30 519
rect 30 -457 64 519
rect -17 -541 17 -507
<< metal1 >>
rect -70 519 -24 531
rect -70 -457 -64 519
rect -30 -457 -24 519
rect -70 -469 -24 -457
rect 24 519 70 531
rect 24 -457 30 519
rect 64 -457 70 519
rect 24 -469 70 -457
rect -29 -507 29 -501
rect -29 -541 -17 -507
rect 17 -541 29 -507
rect -29 -547 29 -541
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.0 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
