* NGSPICE file created from voltage_limiter.ext - technology: sky130A

.subckt voltage_limiter vrec vss vdd
X0 vss.t9 a_4680_n6808.t5 a_3728_n2638.t1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=700000u
X1 a_4680_n6808.t1 a_4680_n6808.t0 a_4750_n2638.t1 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X2 a_3474_n6808.t0 a_4076_n3556.t0 vss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=1.41e+07u
X3 a_4680_n6808.t4 a_4076_n3556.t1 vss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=1.41e+07u
X4 a_7444_n6808.t1 a_8048_n3556.t0 vss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=1.41e+07u
X5 a_8652_n6808.t0 a_8048_n3556.t1 vss.t7 sky130_fd_pr__res_xhigh_po_1p41 l=1.41e+07u
X6 vdd.t15 a_3728_n2638.t2 vss.t13 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X7 a_8652_n6808.t1 vdd.t5 vss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41e+07u
X8 a_4132_n2638.t5 a_4750_n2638.t4 a_4750_n2638.t5 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X9 a_3474_n6808.t1 a_2872_n3556.t1 vss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=1.41e+07u
X10 a_4750_n2638.t3 a_4750_n2638.t2 a_4132_n2638.t4 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X11 vss.t11 a_3728_n2638.t3 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X12 vdd.t11 a_3728_n2638.t4 vss.t12 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X13 vss.t4 a_2872_n3556.t0 vss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41e+07u
X14 vss.t14 a_3728_n2638.t5 vdd.t9 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X15 a_6236_n6808.t0 a_3728_n2638.t0 vss.t6 sky130_fd_pr__res_xhigh_po_1p41 l=1.41e+07u
X16 a_4132_n2638.t3 a_4132_n2638.t2 vdd.t4 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X17 a_6236_n6808.t1 a_6840_n3556.t1 vss.t15 sky130_fd_pr__res_xhigh_po_1p41 l=1.41e+07u
X18 a_4750_n2638.t0 a_4680_n6808.t2 a_4680_n6808.t3 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X19 vdd.t2 a_4132_n2638.t0 a_4132_n2638.t1 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=350000u
X20 a_7444_n6808.t0 a_6840_n3556.t0 vss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41e+07u
X21 vrec.t0 vdd.t0 vss sky130_fd_pr__res_xhigh_po_5p73 l=500000u
R0 a_4680_n6808.n0 a_4680_n6808.t2 319.68
R1 a_4680_n6808.n0 a_4680_n6808.t0 319.675
R2 a_4680_n6808.t5 a_4680_n6808.n1 90.609
R3 a_4680_n6808.t4 a_4680_n6808.t5 89.65
R4 a_4680_n6808.n1 a_4680_n6808.t3 7.141
R5 a_4680_n6808.n1 a_4680_n6808.t1 7.141
R6 a_4680_n6808.n1 a_4680_n6808.n0 0.537
R7 a_3728_n2638.n0 a_3728_n2638.t5 319.852
R8 a_3728_n2638.n0 a_3728_n2638.t4 319.803
R9 a_3728_n2638.n1 a_3728_n2638.t2 159.915
R10 a_3728_n2638.n1 a_3728_n2638.t3 159.892
R11 a_3728_n2638.n2 a_3728_n2638.n1 80.629
R12 a_3728_n2638.t0 a_3728_n2638.t1 12.726
R13 a_3728_n2638.n2 a_3728_n2638.n0 2.831
R14 a_3728_n2638.t0 a_3728_n2638.n2 1.006
R15 vss.n33 vss.t10 397.967
R16 vss.n28 vss.t8 363.009
R17 vss.n31 vss.t15 362.848
R18 vss.n29 vss.t2 362.848
R19 vss.n28 vss.t7 362.848
R20 vss.n25 vss.t6 361.89
R21 vss.n27 vss.t0 361.889
R22 vss.n35 vss.t5 360.459
R23 vss.n37 vss.t3 359.82
R24 vss.n1 vss.t1 359.5
R25 vss.n7 vss.n6 9.3
R26 vss.n10 vss.n9 9.3
R27 vss.n12 vss.n11 9.3
R28 vss.n15 vss.n14 9.3
R29 vss.n22 vss.n21 9.3
R30 vss.n19 vss.n18 9.3
R31 vss.n9 vss.n8 9.154
R32 vss.n14 vss.n13 9.154
R33 vss.n21 vss.n20 9.154
R34 vss.n24 vss.t9 8.704
R35 vss.n0 vss.t12 7.141
R36 vss.n0 vss.t14 7.141
R37 vss.n26 vss.t13 7.141
R38 vss.n26 vss.t11 7.141
R39 vss.n5 vss.n4 6.207
R40 vss.n17 vss.n16 5.949
R41 vss.n3 vss.n2 5.647
R42 vss.n24 vss.n3 3.033
R43 vss.n27 vss.n26 1.732
R44 vss.n1 vss.n0 1.618
R45 vss.n32 vss.n25 0.958
R46 vss.n34 vss.n1 0.956
R47 vss.n30 vss.n27 0.956
R48 vss vss.n37 0.523
R49 vss.n33 vss.n32 0.415
R50 vss.n36 vss.t4 0.351
R51 vss.n25 vss.n24 0.234
R52 vss.n29 vss.n28 0.161
R53 vss.n30 vss.n29 0.161
R54 vss.n31 vss.n30 0.161
R55 vss.n32 vss.n31 0.161
R56 vss.n34 vss.n33 0.16
R57 vss.n35 vss.n34 0.16
R58 vss.n37 vss.n36 0.105
R59 vss.n36 vss.n35 0.08
R60 vss.n19 vss.n17 0.052
R61 vss.n7 vss.n5 0.044
R62 vss.n22 vss.n19 0.035
R63 vss.n23 vss.n22 0.035
R64 vss.n15 vss.n12 0.035
R65 vss.n12 vss.n10 0.035
R66 vss.n10 vss.n7 0.035
R67 vss.n24 vss.n15 0.019
R68 vss.n24 vss.n23 0.015
R69 a_4750_n2638.n1 a_4750_n2638.t4 320.741
R70 a_4750_n2638.n0 a_4750_n2638.t2 320.728
R71 a_4750_n2638.n2 a_4750_n2638.t0 8.198
R72 a_4750_n2638.t1 a_4750_n2638.n3 8.198
R73 a_4750_n2638.n0 a_4750_n2638.t3 7.141
R74 a_4750_n2638.n1 a_4750_n2638.t5 7.141
R75 a_4750_n2638.n3 a_4750_n2638.n0 1.471
R76 a_4750_n2638.n2 a_4750_n2638.n1 1.471
R77 a_4750_n2638.n3 a_4750_n2638.n2 0.331
R78 vdd.n58 vdd.t16 156.029
R79 vdd.n162 vdd.t17 156.029
R80 vdd.n5 vdd.t3 136.278
R81 vdd.n5 vdd.t10 136.278
R82 vdd.n385 vdd.t8 136.278
R83 vdd.n214 vdd.t14 136.278
R84 vdd.n265 vdd.t12 136.278
R85 vdd.n265 vdd.t1 136.278
R86 vdd.n131 vdd.t6 131.1
R87 vdd.n350 vdd.t7 131.1
R88 vdd.n324 vdd.n323 16.607
R89 vdd.n109 vdd.n106 12.969
R90 vdd.n329 vdd.n325 12.968
R91 vdd.n65 vdd.n62 12.745
R92 vdd.n169 vdd.n166 12.745
R93 vdd.n221 vdd.n218 12.698
R94 vdd.n393 vdd.n389 12.697
R95 vdd.n14 vdd.n11 12.685
R96 vdd.n273 vdd.n269 12.685
R97 vdd.n383 vdd.n382 12.369
R98 vdd.n437 vdd.n436 9.3
R99 vdd.n395 vdd.n394 9.3
R100 vdd.n401 vdd.n400 9.3
R101 vdd.n407 vdd.n406 9.3
R102 vdd.n415 vdd.n414 9.3
R103 vdd.n421 vdd.n420 9.3
R104 vdd.n427 vdd.n426 9.3
R105 vdd.n432 vdd.n431 9.3
R106 vdd.n399 vdd.n398 9.3
R107 vdd.n405 vdd.n404 9.3
R108 vdd.n419 vdd.n418 9.3
R109 vdd.n425 vdd.n424 9.3
R110 vdd.n430 vdd.n429 9.3
R111 vdd.n435 vdd.n434 9.3
R112 vdd.n16 vdd.n15 9.3
R113 vdd.n19 vdd.n18 9.3
R114 vdd.n21 vdd.n20 9.3
R115 vdd.n24 vdd.n23 9.3
R116 vdd.n26 vdd.n25 9.3
R117 vdd.n31 vdd.n30 9.3
R118 vdd.n34 vdd.n33 9.3
R119 vdd.n36 vdd.n35 9.3
R120 vdd.n39 vdd.n38 9.3
R121 vdd.n41 vdd.n40 9.3
R122 vdd.n44 vdd.n43 9.3
R123 vdd.n46 vdd.n45 9.3
R124 vdd.n49 vdd.n48 9.3
R125 vdd.n51 vdd.n50 9.3
R126 vdd.n67 vdd.n66 9.3
R127 vdd.n70 vdd.n69 9.3
R128 vdd.n72 vdd.n71 9.3
R129 vdd.n75 vdd.n74 9.3
R130 vdd.n77 vdd.n76 9.3
R131 vdd.n83 vdd.n82 9.3
R132 vdd.n86 vdd.n85 9.3
R133 vdd.n88 vdd.n87 9.3
R134 vdd.n91 vdd.n90 9.3
R135 vdd.n93 vdd.n92 9.3
R136 vdd.n96 vdd.n95 9.3
R137 vdd.n98 vdd.n97 9.3
R138 vdd.n101 vdd.n100 9.3
R139 vdd.n103 vdd.n102 9.3
R140 vdd.n331 vdd.n330 9.3
R141 vdd.n337 vdd.n336 9.3
R142 vdd.n343 vdd.n342 9.3
R143 vdd.n349 vdd.n348 9.3
R144 vdd.n360 vdd.n359 9.3
R145 vdd.n366 vdd.n365 9.3
R146 vdd.n372 vdd.n371 9.3
R147 vdd.n377 vdd.n376 9.3
R148 vdd.n335 vdd.n334 9.3
R149 vdd.n341 vdd.n340 9.3
R150 vdd.n347 vdd.n346 9.3
R151 vdd.n364 vdd.n363 9.3
R152 vdd.n370 vdd.n369 9.3
R153 vdd.n375 vdd.n374 9.3
R154 vdd.n111 vdd.n110 9.3
R155 vdd.n114 vdd.n113 9.3
R156 vdd.n116 vdd.n115 9.3
R157 vdd.n119 vdd.n118 9.3
R158 vdd.n121 vdd.n120 9.3
R159 vdd.n124 vdd.n123 9.3
R160 vdd.n126 vdd.n125 9.3
R161 vdd.n140 vdd.n139 9.3
R162 vdd.n143 vdd.n142 9.3
R163 vdd.n145 vdd.n144 9.3
R164 vdd.n148 vdd.n147 9.3
R165 vdd.n150 vdd.n149 9.3
R166 vdd.n153 vdd.n152 9.3
R167 vdd.n155 vdd.n154 9.3
R168 vdd.n171 vdd.n170 9.3
R169 vdd.n174 vdd.n173 9.3
R170 vdd.n176 vdd.n175 9.3
R171 vdd.n179 vdd.n178 9.3
R172 vdd.n181 vdd.n180 9.3
R173 vdd.n187 vdd.n186 9.3
R174 vdd.n190 vdd.n189 9.3
R175 vdd.n192 vdd.n191 9.3
R176 vdd.n195 vdd.n194 9.3
R177 vdd.n197 vdd.n196 9.3
R178 vdd.n200 vdd.n199 9.3
R179 vdd.n202 vdd.n201 9.3
R180 vdd.n205 vdd.n204 9.3
R181 vdd.n207 vdd.n206 9.3
R182 vdd.n275 vdd.n274 9.3
R183 vdd.n281 vdd.n280 9.3
R184 vdd.n287 vdd.n286 9.3
R185 vdd.n295 vdd.n294 9.3
R186 vdd.n301 vdd.n300 9.3
R187 vdd.n307 vdd.n306 9.3
R188 vdd.n313 vdd.n312 9.3
R189 vdd.n318 vdd.n317 9.3
R190 vdd.n279 vdd.n278 9.3
R191 vdd.n285 vdd.n284 9.3
R192 vdd.n299 vdd.n298 9.3
R193 vdd.n305 vdd.n304 9.3
R194 vdd.n311 vdd.n310 9.3
R195 vdd.n316 vdd.n315 9.3
R196 vdd.n223 vdd.n222 9.3
R197 vdd.n226 vdd.n225 9.3
R198 vdd.n228 vdd.n227 9.3
R199 vdd.n231 vdd.n230 9.3
R200 vdd.n233 vdd.n232 9.3
R201 vdd.n240 vdd.n239 9.3
R202 vdd.n243 vdd.n242 9.3
R203 vdd.n245 vdd.n244 9.3
R204 vdd.n248 vdd.n247 9.3
R205 vdd.n250 vdd.n249 9.3
R206 vdd.n253 vdd.n252 9.3
R207 vdd.n255 vdd.n254 9.3
R208 vdd.n258 vdd.n257 9.3
R209 vdd.n260 vdd.n259 9.3
R210 vdd.n392 vdd.n391 8.855
R211 vdd.n398 vdd.n397 8.855
R212 vdd.n404 vdd.n403 8.855
R213 vdd.n410 vdd.n409 8.855
R214 vdd.n388 vdd.n387 8.855
R215 vdd.n418 vdd.n417 8.855
R216 vdd.n424 vdd.n423 8.855
R217 vdd.n429 vdd.n428 8.855
R218 vdd.n434 vdd.n433 8.855
R219 vdd.n13 vdd.n12 8.855
R220 vdd.n18 vdd.n17 8.855
R221 vdd.n23 vdd.n22 8.855
R222 vdd.n10 vdd.n9 8.855
R223 vdd.n8 vdd.n7 8.855
R224 vdd.n33 vdd.n32 8.855
R225 vdd.n38 vdd.n37 8.855
R226 vdd.n43 vdd.n42 8.855
R227 vdd.n48 vdd.n47 8.855
R228 vdd.n64 vdd.n63 8.855
R229 vdd.n69 vdd.n68 8.855
R230 vdd.n74 vdd.n73 8.855
R231 vdd.n79 vdd.n78 8.855
R232 vdd.n61 vdd.n60 8.855
R233 vdd.n85 vdd.n84 8.855
R234 vdd.n90 vdd.n89 8.855
R235 vdd.n95 vdd.n94 8.855
R236 vdd.n100 vdd.n99 8.855
R237 vdd.n328 vdd.n327 8.855
R238 vdd.n334 vdd.n333 8.855
R239 vdd.n340 vdd.n339 8.855
R240 vdd.n346 vdd.n345 8.855
R241 vdd.n353 vdd.n352 8.855
R242 vdd.n357 vdd.n356 8.855
R243 vdd.n363 vdd.n362 8.855
R244 vdd.n369 vdd.n368 8.855
R245 vdd.n374 vdd.n373 8.855
R246 vdd.n108 vdd.n107 8.855
R247 vdd.n113 vdd.n112 8.855
R248 vdd.n118 vdd.n117 8.855
R249 vdd.n123 vdd.n122 8.855
R250 vdd.n134 vdd.n133 8.855
R251 vdd.n137 vdd.n136 8.855
R252 vdd.n142 vdd.n141 8.855
R253 vdd.n147 vdd.n146 8.855
R254 vdd.n152 vdd.n151 8.855
R255 vdd.n168 vdd.n167 8.855
R256 vdd.n173 vdd.n172 8.855
R257 vdd.n178 vdd.n177 8.855
R258 vdd.n183 vdd.n182 8.855
R259 vdd.n165 vdd.n164 8.855
R260 vdd.n189 vdd.n188 8.855
R261 vdd.n194 vdd.n193 8.855
R262 vdd.n199 vdd.n198 8.855
R263 vdd.n204 vdd.n203 8.855
R264 vdd.n272 vdd.n271 8.855
R265 vdd.n278 vdd.n277 8.855
R266 vdd.n284 vdd.n283 8.855
R267 vdd.n290 vdd.n289 8.855
R268 vdd.n268 vdd.n267 8.855
R269 vdd.n298 vdd.n297 8.855
R270 vdd.n304 vdd.n303 8.855
R271 vdd.n310 vdd.n309 8.855
R272 vdd.n315 vdd.n314 8.855
R273 vdd.n220 vdd.n219 8.855
R274 vdd.n225 vdd.n224 8.855
R275 vdd.n230 vdd.n229 8.855
R276 vdd.n235 vdd.n234 8.855
R277 vdd.n217 vdd.n216 8.855
R278 vdd.n242 vdd.n241 8.855
R279 vdd.n247 vdd.n246 8.855
R280 vdd.n252 vdd.n251 8.855
R281 vdd.n257 vdd.n256 8.855
R282 vdd.n133 vdd.n132 7.775
R283 vdd.n216 vdd.n215 7.775
R284 vdd.n60 vdd.n59 7.49
R285 vdd.n164 vdd.n163 7.49
R286 vdd.n7 vdd.n6 7.463
R287 vdd.n28 vdd.t4 7.141
R288 vdd.n412 vdd.t9 7.141
R289 vdd.n28 vdd.t11 7.141
R290 vdd.n292 vdd.t13 7.141
R291 vdd.n292 vdd.t2 7.141
R292 vdd.n237 vdd.t15 7.141
R293 vdd.n52 vdd.n0 6.209
R294 vdd.n319 vdd.n263 6.209
R295 vdd.n438 vdd.n383 6.207
R296 vdd.n261 vdd.n209 6.207
R297 vdd.n104 vdd.n53 6.201
R298 vdd.n208 vdd.n157 6.201
R299 vdd.n27 vdd.n10 5.985
R300 vdd.n291 vdd.n290 5.985
R301 vdd.n411 vdd.n410 5.982
R302 vdd.n236 vdd.n235 5.982
R303 vdd.n80 vdd.n79 5.969
R304 vdd.n358 vdd.n357 5.969
R305 vdd.n138 vdd.n137 5.969
R306 vdd.n184 vdd.n183 5.969
R307 vdd.n266 vdd.n265 5.95
R308 vdd.n378 vdd.n324 5.735
R309 vdd.n156 vdd.n105 5.735
R310 vdd.n273 vdd.n272 5.606
R311 vdd.n14 vdd.n13 5.606
R312 vdd.n393 vdd.n392 5.603
R313 vdd.n221 vdd.n220 5.603
R314 vdd.n65 vdd.n64 5.592
R315 vdd.n169 vdd.n168 5.592
R316 vdd.n329 vdd.n328 5.56
R317 vdd.n109 vdd.n108 5.56
R318 vdd.n386 vdd.n385 5.347
R319 vdd.n351 vdd.n350 5.347
R320 vdd.n423 vdd.n422 3.685
R321 vdd.n417 vdd.n416 3.685
R322 vdd.n387 vdd.n386 3.685
R323 vdd.n409 vdd.n408 3.685
R324 vdd.n403 vdd.n402 3.685
R325 vdd.n397 vdd.n396 3.685
R326 vdd.n368 vdd.n367 3.685
R327 vdd.n362 vdd.n361 3.685
R328 vdd.n356 vdd.n355 3.685
R329 vdd.n352 vdd.n351 3.685
R330 vdd.n345 vdd.n344 3.685
R331 vdd.n339 vdd.n338 3.685
R332 vdd.n333 vdd.n332 3.685
R333 vdd.n391 vdd.n390 3.514
R334 vdd.n327 vdd.n326 3.514
R335 vdd.n29 vdd.n8 3.512
R336 vdd.n293 vdd.n268 3.512
R337 vdd.n413 vdd.n388 3.511
R338 vdd.n238 vdd.n217 3.511
R339 vdd.n81 vdd.n61 3.507
R340 vdd.n354 vdd.n353 3.507
R341 vdd.n135 vdd.n134 3.507
R342 vdd.n185 vdd.n165 3.507
R343 vdd.n309 vdd.n308 3.052
R344 vdd.n303 vdd.n302 3.052
R345 vdd.n297 vdd.n296 3.052
R346 vdd.n267 vdd.n266 3.052
R347 vdd.n289 vdd.n288 3.052
R348 vdd.n283 vdd.n282 3.052
R349 vdd.n277 vdd.n276 3.052
R350 vdd.n271 vdd.n270 2.91
R351 vdd.n440 vdd.t0 2.699
R352 vdd.n262 vdd.t5 1.64
R353 vdd.n379 vdd.n378 1.601
R354 vdd.n322 vdd.n156 1.601
R355 vdd.n380 vdd.n104 1.551
R356 vdd.n321 vdd.n208 1.551
R357 vdd.n439 vdd.n438 0.798
R358 vdd.n262 vdd.n261 0.798
R359 vdd.n381 vdd.n52 0.785
R360 vdd.n320 vdd.n319 0.785
R361 vdd.n111 vdd.n109 0.772
R362 vdd.n331 vdd.n329 0.772
R363 vdd.n67 vdd.n65 0.735
R364 vdd.n171 vdd.n169 0.735
R365 vdd.n265 vdd.n264 0.729
R366 vdd.n5 vdd.n4 0.697
R367 vdd.n5 vdd.n3 0.697
R368 vdd.n6 vdd.n5 0.697
R369 vdd.n5 vdd.n2 0.697
R370 vdd.n5 vdd.n1 0.697
R371 vdd.n58 vdd.n57 0.683
R372 vdd.n58 vdd.n56 0.683
R373 vdd.n59 vdd.n58 0.683
R374 vdd.n58 vdd.n55 0.683
R375 vdd.n58 vdd.n54 0.683
R376 vdd.n162 vdd.n161 0.683
R377 vdd.n162 vdd.n160 0.683
R378 vdd.n163 vdd.n162 0.683
R379 vdd.n162 vdd.n159 0.683
R380 vdd.n162 vdd.n158 0.683
R381 vdd.n223 vdd.n221 0.677
R382 vdd.n395 vdd.n393 0.677
R383 vdd.n16 vdd.n14 0.662
R384 vdd.n275 vdd.n273 0.662
R385 vdd.n385 vdd.n384 0.592
R386 vdd.n131 vdd.n130 0.54
R387 vdd.n131 vdd.n129 0.54
R388 vdd.n132 vdd.n131 0.54
R389 vdd.n131 vdd.n128 0.54
R390 vdd.n131 vdd.n127 0.54
R391 vdd.n214 vdd.n213 0.54
R392 vdd.n214 vdd.n212 0.54
R393 vdd.n215 vdd.n214 0.54
R394 vdd.n214 vdd.n211 0.54
R395 vdd.n214 vdd.n210 0.54
R396 vdd.n440 vdd.n439 0.497
R397 vdd vdd.n440 0.301
R398 vdd.n322 vdd.n321 0.159
R399 vdd.n380 vdd.n379 0.159
R400 vdd.n321 vdd.n320 0.151
R401 vdd.n381 vdd.n380 0.151
R402 vdd.n379 vdd.n322 0.111
R403 vdd.n80 vdd.n77 0.108
R404 vdd.n360 vdd.n358 0.108
R405 vdd.n140 vdd.n138 0.108
R406 vdd.n184 vdd.n181 0.108
R407 vdd.n320 vdd.n262 0.107
R408 vdd.n439 vdd.n381 0.107
R409 vdd.n378 vdd.n377 0.106
R410 vdd.n156 vdd.n155 0.106
R411 vdd.n83 vdd.n81 0.093
R412 vdd.n354 vdd.n349 0.093
R413 vdd.n135 vdd.n126 0.093
R414 vdd.n187 vdd.n185 0.093
R415 vdd.n81 vdd.n80 0.093
R416 vdd.n358 vdd.n354 0.093
R417 vdd.n138 vdd.n135 0.093
R418 vdd.n185 vdd.n184 0.093
R419 vdd.n104 vdd.n103 0.091
R420 vdd.n208 vdd.n207 0.091
R421 vdd.n103 vdd.n101 0.073
R422 vdd.n101 vdd.n98 0.073
R423 vdd.n98 vdd.n96 0.073
R424 vdd.n96 vdd.n93 0.073
R425 vdd.n93 vdd.n91 0.073
R426 vdd.n91 vdd.n88 0.073
R427 vdd.n88 vdd.n86 0.073
R428 vdd.n86 vdd.n83 0.073
R429 vdd.n77 vdd.n75 0.073
R430 vdd.n75 vdd.n72 0.073
R431 vdd.n72 vdd.n70 0.073
R432 vdd.n70 vdd.n67 0.073
R433 vdd.n377 vdd.n375 0.073
R434 vdd.n375 vdd.n372 0.073
R435 vdd.n372 vdd.n370 0.073
R436 vdd.n370 vdd.n366 0.073
R437 vdd.n366 vdd.n364 0.073
R438 vdd.n364 vdd.n360 0.073
R439 vdd.n349 vdd.n347 0.073
R440 vdd.n347 vdd.n343 0.073
R441 vdd.n343 vdd.n341 0.073
R442 vdd.n341 vdd.n337 0.073
R443 vdd.n337 vdd.n335 0.073
R444 vdd.n335 vdd.n331 0.073
R445 vdd.n155 vdd.n153 0.073
R446 vdd.n153 vdd.n150 0.073
R447 vdd.n150 vdd.n148 0.073
R448 vdd.n148 vdd.n145 0.073
R449 vdd.n145 vdd.n143 0.073
R450 vdd.n143 vdd.n140 0.073
R451 vdd.n126 vdd.n124 0.073
R452 vdd.n124 vdd.n121 0.073
R453 vdd.n121 vdd.n119 0.073
R454 vdd.n119 vdd.n116 0.073
R455 vdd.n116 vdd.n114 0.073
R456 vdd.n114 vdd.n111 0.073
R457 vdd.n207 vdd.n205 0.073
R458 vdd.n205 vdd.n202 0.073
R459 vdd.n202 vdd.n200 0.073
R460 vdd.n200 vdd.n197 0.073
R461 vdd.n197 vdd.n195 0.073
R462 vdd.n195 vdd.n192 0.073
R463 vdd.n192 vdd.n190 0.073
R464 vdd.n190 vdd.n187 0.073
R465 vdd.n181 vdd.n179 0.073
R466 vdd.n179 vdd.n176 0.073
R467 vdd.n176 vdd.n174 0.073
R468 vdd.n174 vdd.n171 0.073
R469 vdd.n411 vdd.n407 0.048
R470 vdd.n236 vdd.n233 0.048
R471 vdd.n415 vdd.n413 0.041
R472 vdd.n240 vdd.n238 0.041
R473 vdd.n438 vdd.n437 0.04
R474 vdd.n261 vdd.n260 0.04
R475 vdd.n412 vdd.n411 0.036
R476 vdd.n237 vdd.n236 0.036
R477 vdd.n437 vdd.n435 0.032
R478 vdd.n435 vdd.n432 0.032
R479 vdd.n432 vdd.n430 0.032
R480 vdd.n430 vdd.n427 0.032
R481 vdd.n427 vdd.n425 0.032
R482 vdd.n425 vdd.n421 0.032
R483 vdd.n421 vdd.n419 0.032
R484 vdd.n419 vdd.n415 0.032
R485 vdd.n407 vdd.n405 0.032
R486 vdd.n405 vdd.n401 0.032
R487 vdd.n401 vdd.n399 0.032
R488 vdd.n399 vdd.n395 0.032
R489 vdd.n260 vdd.n258 0.032
R490 vdd.n258 vdd.n255 0.032
R491 vdd.n255 vdd.n253 0.032
R492 vdd.n253 vdd.n250 0.032
R493 vdd.n250 vdd.n248 0.032
R494 vdd.n248 vdd.n245 0.032
R495 vdd.n245 vdd.n243 0.032
R496 vdd.n243 vdd.n240 0.032
R497 vdd.n233 vdd.n231 0.032
R498 vdd.n231 vdd.n228 0.032
R499 vdd.n228 vdd.n226 0.032
R500 vdd.n226 vdd.n223 0.032
R501 vdd.n27 vdd.n26 0.032
R502 vdd.n291 vdd.n287 0.032
R503 vdd.n31 vdd.n29 0.027
R504 vdd.n295 vdd.n293 0.027
R505 vdd.n52 vdd.n51 0.027
R506 vdd.n319 vdd.n318 0.027
R507 vdd.n28 vdd.n27 0.024
R508 vdd.n292 vdd.n291 0.024
R509 vdd.n51 vdd.n49 0.021
R510 vdd.n49 vdd.n46 0.021
R511 vdd.n46 vdd.n44 0.021
R512 vdd.n44 vdd.n41 0.021
R513 vdd.n41 vdd.n39 0.021
R514 vdd.n39 vdd.n36 0.021
R515 vdd.n36 vdd.n34 0.021
R516 vdd.n34 vdd.n31 0.021
R517 vdd.n26 vdd.n24 0.021
R518 vdd.n24 vdd.n21 0.021
R519 vdd.n21 vdd.n19 0.021
R520 vdd.n19 vdd.n16 0.021
R521 vdd.n318 vdd.n316 0.021
R522 vdd.n316 vdd.n313 0.021
R523 vdd.n313 vdd.n311 0.021
R524 vdd.n311 vdd.n307 0.021
R525 vdd.n307 vdd.n305 0.021
R526 vdd.n305 vdd.n301 0.021
R527 vdd.n301 vdd.n299 0.021
R528 vdd.n299 vdd.n295 0.021
R529 vdd.n287 vdd.n285 0.021
R530 vdd.n285 vdd.n281 0.021
R531 vdd.n281 vdd.n279 0.021
R532 vdd.n279 vdd.n275 0.021
R533 vdd.n413 vdd.n412 0.006
R534 vdd.n238 vdd.n237 0.006
R535 vdd.n29 vdd.n28 0.004
R536 vdd.n293 vdd.n292 0.004
R537 a_3474_n6808.t0 a_3474_n6808.t1 0.179
R538 a_4076_n3556.t0 a_4076_n3556.t1 0.179
R539 a_7444_n6808.t0 a_7444_n6808.t1 0.179
R540 a_8048_n3556.t0 a_8048_n3556.t1 0.179
R541 a_8652_n6808.t0 a_8652_n6808.t1 0.179
R542 a_4132_n2638.n0 a_4132_n2638.t0 320.353
R543 a_4132_n2638.n3 a_4132_n2638.t2 320.262
R544 a_4132_n2638.n1 a_4132_n2638.t5 8.177
R545 a_4132_n2638.n2 a_4132_n2638.t4 7.978
R546 a_4132_n2638.n0 a_4132_n2638.t1 7.141
R547 a_4132_n2638.t3 a_4132_n2638.n3 7.141
R548 a_4132_n2638.n2 a_4132_n2638.n1 1.561
R549 a_4132_n2638.n1 a_4132_n2638.n0 1.351
R550 a_4132_n2638.n3 a_4132_n2638.n2 1.261
R551 a_2872_n3556.t0 a_2872_n3556.t1 0.179
R552 a_6236_n6808.t0 a_6236_n6808.t1 0.179
R553 a_6840_n3556.t0 a_6840_n3556.t1 0.179
R554 vrec.n0 vrec.t0 2.413
R555 vrec vrec.n0 0.248
R556 vrec.n0 vrec 0.069
C0 vrec vdd 1.58fF
.ends

