* NGSPICE file created from Temperature_Sensor.ext - technology: sky130A

.subckt Temperature_Sensor vtemp vss vdd
X0 a_n3070_n3662.t10 a_n3836_n1894.t3 vdd.t27 vss.t20 sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=8.6 as=0.58 ps=4.29 w=4 l=2
X1 a_n3070_n3662.t9 a_n3836_n1894.t4 vdd.t22 vss.t17 sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=8.6 as=0.58 ps=4.29 w=4 l=2
X2 a_n5752_n3086# a_n5752_n2774# a_n5810_n2748# vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=0.6 pd=4.6 as=0.58 ps=4.58 w=2 l=2
X3 a_n178_n2405.t10 a_n178_n2405.t9 vdd.t9 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=1.5 ps=10.6 w=5 l=2
X4 a_n3216_n2108.t0 a_n3836_n1894.t1 a_n3836_n1894.t2 vss.t21 sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=8.6 as=1.16 ps=8.58 w=4 l=2
X5 vdd.t3 a_n178_n2405.t7 a_n178_n2405.t8 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X6 vdd.t20 a_n3836_n1894.t5 a_n3070_n3662.t8 vss.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.2 ps=8.6 w=4 l=2
X7 a_n178_n2405.t6 a_n178_n2405.t5 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=1.5 ps=10.6 w=5 l=2
X8 vss.t16 a_n5752_n2774# a_n5752_n2774# vss.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.15 ps=1.6 w=0.5 l=2
X9 vtemp.t3 a_n3070_n3662.t11 a_62_n3136# vss.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.3 ps=2.6 w=1 l=0.5
X10 a_62_n3136# a_n3216_n2108.t2 a_n178_n2405.t1 vss.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.145 ps=1.29 w=1 l=2
X11 vdd.t26 a_n3836_n1894.t6 a_n3070_n3662.t7 vss.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.2 ps=8.6 w=4 l=2
X12 vss.t14 a_n5752_n2774# a_62_n3136# vss.t13 sky130_fd_pr__nfet_01v8 ad=1.5 pd=10.6 as=1.45 ps=10.6 w=5 l=2
X13 vss.t12 a_n5752_n2774# a_62_n3136# vss.t11 sky130_fd_pr__nfet_01v8 ad=1.5 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X14 vss.t28 vss.t27 a_n3216_n2108.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
X15 a_n5752_n1958# a_n5752_n1958# vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.6 ps=4.6 w=2 l=2
X16 vdd.t24 a_n3836_n1894.t7 a_n3070_n3662.t6 vss.t17 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.2 ps=8.6 w=4 l=2
X17 a_n3070_n3662.t5 a_n3836_n1894.t8 vdd.t25 vss.t20 sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=8.6 as=0.58 ps=4.29 w=4 l=2
X18 vss.t26 vss.t25 a_n3070_n3662.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
X19 a_62_n3136# a_n3216_n2108.t3 a_n178_n2405.t2 vss.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.145 ps=1.29 w=1 l=2
X20 a_62_n3136# a_n5752_n2774# vss.t10 vss.t9 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.5 ps=10.6 w=5 l=2
X21 vdd.t5 a_n178_n2405.t12 vtemp.t7 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X22 vtemp.t6 a_n178_n2405.t13 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=1.5 ps=10.6 w=5 l=2
X23 vtemp.t2 a_n3070_n3662.t12 a_62_n3136# vss.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.3 ps=2.6 w=1 l=0.5
X24 a_n178_n2405.t11 a_n3216_n2108.t4 a_62_n3136# vss.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.3 ps=2.6 w=1 l=2
X25 a_n178_n2405.t0 a_n3216_n2108.t5 a_62_n3136# vss.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.3 ps=2.6 w=1 l=2
X26 a_n3070_n3662.t4 a_n3836_n1894.t9 vdd.t29 vss.t17 sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=8.6 as=0.58 ps=4.29 w=4 l=2
X27 a_n3836_n1894.t0 a_n5752_n2774# vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.6 ps=4.6 w=2 l=2
X28 a_n5752_n1958# a_n5752_n2774# a_n5752_n2774# vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.6 ps=4.6 w=2 l=2
X29 a_n5752_n3086# a_n5752_n3086# vss.t23 vss.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.145 ps=1.58 w=0.5 l=2
X30 a_62_n3136# a_n3070_n3662.t13 vtemp.t1 vss.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.145 ps=1.29 w=1 l=0.5
X31 vdd.t28 a_n3836_n1894.t10 a_n3070_n3662.t3 vss.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.2 ps=8.6 w=4 l=2
X32 vdd.t23 a_n3836_n1894.t11 a_n3070_n3662.t2 vss.t18 sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.2 ps=8.6 w=4 l=2
X33 vdd.t13 a_n5752_n1958# a_n5810_n2748# vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=0.6 pd=4.6 as=0.58 ps=4.58 w=2 l=2
X34 vtemp.t5 a_n178_n2405.t14 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=1.5 ps=10.6 w=5 l=2
X35 a_62_n3136# a_n5752_n2774# vss.t8 vss.t7 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.5 ps=10.6 w=5 l=2
X36 vdd.t31 a_n178_n2405.t15 vtemp.t4 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X37 vdd.t7 a_n178_n2405.t3 a_n178_n2405.t4 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X38 a_62_n3136# a_n3070_n3662.t14 vtemp.t0 vss.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.145 ps=1.29 w=1 l=0.5
X39 vdd.t21 a_n3836_n1894.t12 a_n3070_n3662.t1 vss.t17 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.2 ps=8.6 w=4 l=2
R0 a_n3836_n1894.n4 a_n3836_n1894.t12 54.8313
R1 a_n3836_n1894.n1 a_n3836_n1894.t9 54.8313
R2 a_n3836_n1894.n2 a_n3836_n1894.t11 54.8313
R3 a_n3836_n1894.n0 a_n3836_n1894.t3 54.8313
R4 a_n3836_n1894.n0 a_n3836_n1894.t8 54.8309
R5 a_n3836_n1894.n1 a_n3836_n1894.t4 54.8309
R6 a_n3836_n1894.n3 a_n3836_n1894.t6 54.8306
R7 a_n3836_n1894.n3 a_n3836_n1894.t10 54.8306
R8 a_n3836_n1894.n2 a_n3836_n1894.t5 54.8306
R9 a_n3836_n1894.n4 a_n3836_n1894.t7 54.8306
R10 a_n3836_n1894.n8 a_n3836_n1894.t1 54.8305
R11 a_n3836_n1894.n9 a_n3836_n1894.t0 14.3139
R12 a_n3836_n1894.t2 a_n3836_n1894.n9 4.35262
R13 a_n3836_n1894.n1 a_n3836_n1894.n4 1.48142
R14 a_n3836_n1894.n9 a_n3836_n1894.n8 1.41958
R15 a_n3836_n1894.n2 a_n3836_n1894.n1 1.3917
R16 a_n3836_n1894.n3 a_n3836_n1894.n0 1.39134
R17 a_n3836_n1894.n8 a_n3836_n1894.n3 1.26382
R18 a_n3836_n1894.n7 a_n3836_n1894.n6 1.263
R19 a_n3836_n1894.n0 a_n3836_n1894.n2 1.263
R20 a_n3836_n1894.n3 a_n3836_n1894.n7 0.955675
R21 a_n3836_n1894.n6 a_n3836_n1894.n5 0.954667
R22 vdd.n422 vdd.t14 512.189
R23 vdd.n422 vdd.t12 512.189
R24 vdd.n427 vdd.t16 512.189
R25 vdd.n427 vdd.t19 512.189
R26 vdd.n400 vdd.t17 512.189
R27 vdd.n7 vdd.t6 247.72
R28 vdd.n72 vdd.t8 247.72
R29 vdd.n72 vdd.t30 247.72
R30 vdd.n151 vdd.t10 247.72
R31 vdd.n151 vdd.t2 247.72
R32 vdd.n230 vdd.t32 247.72
R33 vdd.n230 vdd.t4 247.72
R34 vdd.n309 vdd.t0 247.72
R35 vdd.n11 vdd.n8 20.6743
R36 vdd.n399 vdd.n398 16.6308
R37 vdd.n1 vdd.n0 16.6013
R38 vdd.n311 vdd.n310 16.5774
R39 vdd.n424 vdd.n423 16.318
R40 vdd.n426 vdd.n425 16.318
R41 vdd.n74 vdd.n73 16.289
R42 vdd.n153 vdd.n152 16.289
R43 vdd.n232 vdd.n231 16.289
R44 vdd.n462 vdd.t13 14.2849
R45 vdd.n462 vdd.t15 14.2849
R46 vdd.n413 vdd.t18 14.2849
R47 vdd.n405 vdd.n401 12.9284
R48 vdd.n316 vdd.n312 12.9279
R49 vdd.n237 vdd.n233 12.9133
R50 vdd.n158 vdd.n154 12.9133
R51 vdd.n79 vdd.n75 12.9133
R52 vdd.n432 vdd.n428 12.8695
R53 vdd.n441 vdd.n440 9.3005
R54 vdd.n444 vdd.n443 9.3005
R55 vdd.n446 vdd.n445 9.3005
R56 vdd.n452 vdd.n451 9.3005
R57 vdd.n455 vdd.n454 9.3005
R58 vdd.n465 vdd.n464 9.3005
R59 vdd.n468 vdd.n467 9.3005
R60 vdd.n470 vdd.n469 9.3005
R61 vdd.n407 vdd.n406 9.3005
R62 vdd.n417 vdd.n416 9.3005
R63 vdd.n419 vdd.n418 9.3005
R64 vdd.n318 vdd.n317 9.3005
R65 vdd.n324 vdd.n323 9.3005
R66 vdd.n330 vdd.n329 9.3005
R67 vdd.n336 vdd.n335 9.3005
R68 vdd.n342 vdd.n341 9.3005
R69 vdd.n356 vdd.n355 9.3005
R70 vdd.n362 vdd.n361 9.3005
R71 vdd.n368 vdd.n367 9.3005
R72 vdd.n374 vdd.n373 9.3005
R73 vdd.n380 vdd.n379 9.3005
R74 vdd.n385 vdd.n384 9.3005
R75 vdd.n239 vdd.n238 9.3005
R76 vdd.n245 vdd.n244 9.3005
R77 vdd.n251 vdd.n250 9.3005
R78 vdd.n257 vdd.n256 9.3005
R79 vdd.n263 vdd.n262 9.3005
R80 vdd.n277 vdd.n276 9.3005
R81 vdd.n283 vdd.n282 9.3005
R82 vdd.n289 vdd.n288 9.3005
R83 vdd.n295 vdd.n294 9.3005
R84 vdd.n301 vdd.n300 9.3005
R85 vdd.n306 vdd.n305 9.3005
R86 vdd.n160 vdd.n159 9.3005
R87 vdd.n166 vdd.n165 9.3005
R88 vdd.n172 vdd.n171 9.3005
R89 vdd.n178 vdd.n177 9.3005
R90 vdd.n184 vdd.n183 9.3005
R91 vdd.n198 vdd.n197 9.3005
R92 vdd.n204 vdd.n203 9.3005
R93 vdd.n210 vdd.n209 9.3005
R94 vdd.n216 vdd.n215 9.3005
R95 vdd.n222 vdd.n221 9.3005
R96 vdd.n227 vdd.n226 9.3005
R97 vdd.n81 vdd.n80 9.3005
R98 vdd.n87 vdd.n86 9.3005
R99 vdd.n93 vdd.n92 9.3005
R100 vdd.n99 vdd.n98 9.3005
R101 vdd.n105 vdd.n104 9.3005
R102 vdd.n119 vdd.n118 9.3005
R103 vdd.n125 vdd.n124 9.3005
R104 vdd.n131 vdd.n130 9.3005
R105 vdd.n137 vdd.n136 9.3005
R106 vdd.n143 vdd.n142 9.3005
R107 vdd.n148 vdd.n147 9.3005
R108 vdd.n85 vdd.n84 9.3005
R109 vdd.n91 vdd.n90 9.3005
R110 vdd.n97 vdd.n96 9.3005
R111 vdd.n103 vdd.n102 9.3005
R112 vdd.n109 vdd.n108 9.3005
R113 vdd.n123 vdd.n122 9.3005
R114 vdd.n129 vdd.n128 9.3005
R115 vdd.n135 vdd.n134 9.3005
R116 vdd.n141 vdd.n140 9.3005
R117 vdd.n146 vdd.n145 9.3005
R118 vdd.n164 vdd.n163 9.3005
R119 vdd.n170 vdd.n169 9.3005
R120 vdd.n176 vdd.n175 9.3005
R121 vdd.n182 vdd.n181 9.3005
R122 vdd.n188 vdd.n187 9.3005
R123 vdd.n202 vdd.n201 9.3005
R124 vdd.n208 vdd.n207 9.3005
R125 vdd.n214 vdd.n213 9.3005
R126 vdd.n220 vdd.n219 9.3005
R127 vdd.n225 vdd.n224 9.3005
R128 vdd.n243 vdd.n242 9.3005
R129 vdd.n249 vdd.n248 9.3005
R130 vdd.n255 vdd.n254 9.3005
R131 vdd.n261 vdd.n260 9.3005
R132 vdd.n267 vdd.n266 9.3005
R133 vdd.n281 vdd.n280 9.3005
R134 vdd.n287 vdd.n286 9.3005
R135 vdd.n293 vdd.n292 9.3005
R136 vdd.n299 vdd.n298 9.3005
R137 vdd.n304 vdd.n303 9.3005
R138 vdd.n322 vdd.n321 9.3005
R139 vdd.n328 vdd.n327 9.3005
R140 vdd.n334 vdd.n333 9.3005
R141 vdd.n340 vdd.n339 9.3005
R142 vdd.n346 vdd.n345 9.3005
R143 vdd.n360 vdd.n359 9.3005
R144 vdd.n366 vdd.n365 9.3005
R145 vdd.n372 vdd.n371 9.3005
R146 vdd.n378 vdd.n377 9.3005
R147 vdd.n383 vdd.n382 9.3005
R148 vdd.n13 vdd.n12 9.3005
R149 vdd.n16 vdd.n15 9.3005
R150 vdd.n18 vdd.n17 9.3005
R151 vdd.n21 vdd.n20 9.3005
R152 vdd.n23 vdd.n22 9.3005
R153 vdd.n26 vdd.n25 9.3005
R154 vdd.n28 vdd.n27 9.3005
R155 vdd.n31 vdd.n30 9.3005
R156 vdd.n33 vdd.n32 9.3005
R157 vdd.n36 vdd.n35 9.3005
R158 vdd.n45 vdd.n44 9.3005
R159 vdd.n48 vdd.n47 9.3005
R160 vdd.n50 vdd.n49 9.3005
R161 vdd.n53 vdd.n52 9.3005
R162 vdd.n55 vdd.n54 9.3005
R163 vdd.n58 vdd.n57 9.3005
R164 vdd.n60 vdd.n59 9.3005
R165 vdd.n63 vdd.n62 9.3005
R166 vdd.n65 vdd.n64 9.3005
R167 vdd.n68 vdd.n67 9.3005
R168 vdd.n70 vdd.n69 9.3005
R169 vdd.n454 vdd.n453 8.85536
R170 vdd.n431 vdd.n430 8.85536
R171 vdd.n428 vdd.n427 8.85536
R172 vdd.n435 vdd.n434 8.85536
R173 vdd.n443 vdd.n442 8.85536
R174 vdd.n459 vdd.n458 8.85536
R175 vdd.n467 vdd.n466 8.85536
R176 vdd.n449 vdd.n448 8.85536
R177 vdd.n404 vdd.n403 8.85536
R178 vdd.n401 vdd.n400 8.85536
R179 vdd.n411 vdd.n410 8.85536
R180 vdd.n416 vdd.n415 8.85536
R181 vdd.n78 vdd.n77 8.85536
R182 vdd.n84 vdd.n83 8.85536
R183 vdd.n90 vdd.n89 8.85536
R184 vdd.n96 vdd.n95 8.85536
R185 vdd.n102 vdd.n101 8.85536
R186 vdd.n108 vdd.n107 8.85536
R187 vdd.n113 vdd.n112 8.85536
R188 vdd.n122 vdd.n121 8.85536
R189 vdd.n128 vdd.n127 8.85536
R190 vdd.n134 vdd.n133 8.85536
R191 vdd.n140 vdd.n139 8.85536
R192 vdd.n145 vdd.n144 8.85536
R193 vdd.n157 vdd.n156 8.85536
R194 vdd.n163 vdd.n162 8.85536
R195 vdd.n169 vdd.n168 8.85536
R196 vdd.n175 vdd.n174 8.85536
R197 vdd.n181 vdd.n180 8.85536
R198 vdd.n187 vdd.n186 8.85536
R199 vdd.n192 vdd.n191 8.85536
R200 vdd.n201 vdd.n200 8.85536
R201 vdd.n207 vdd.n206 8.85536
R202 vdd.n213 vdd.n212 8.85536
R203 vdd.n219 vdd.n218 8.85536
R204 vdd.n224 vdd.n223 8.85536
R205 vdd.n236 vdd.n235 8.85536
R206 vdd.n242 vdd.n241 8.85536
R207 vdd.n248 vdd.n247 8.85536
R208 vdd.n254 vdd.n253 8.85536
R209 vdd.n260 vdd.n259 8.85536
R210 vdd.n266 vdd.n265 8.85536
R211 vdd.n271 vdd.n270 8.85536
R212 vdd.n280 vdd.n279 8.85536
R213 vdd.n286 vdd.n285 8.85536
R214 vdd.n292 vdd.n291 8.85536
R215 vdd.n298 vdd.n297 8.85536
R216 vdd.n303 vdd.n302 8.85536
R217 vdd.n315 vdd.n314 8.85536
R218 vdd.n321 vdd.n320 8.85536
R219 vdd.n327 vdd.n326 8.85536
R220 vdd.n333 vdd.n332 8.85536
R221 vdd.n339 vdd.n338 8.85536
R222 vdd.n345 vdd.n344 8.85536
R223 vdd.n350 vdd.n349 8.85536
R224 vdd.n359 vdd.n358 8.85536
R225 vdd.n365 vdd.n364 8.85536
R226 vdd.n371 vdd.n370 8.85536
R227 vdd.n377 vdd.n376 8.85536
R228 vdd.n382 vdd.n381 8.85536
R229 vdd.n10 vdd.n9 8.85536
R230 vdd.n15 vdd.n14 8.85536
R231 vdd.n20 vdd.n19 8.85536
R232 vdd.n25 vdd.n24 8.85536
R233 vdd.n30 vdd.n29 8.85536
R234 vdd.n35 vdd.n34 8.85536
R235 vdd.n39 vdd.n38 8.85536
R236 vdd.n47 vdd.n46 8.85536
R237 vdd.n52 vdd.n51 8.85536
R238 vdd.n57 vdd.n56 8.85536
R239 vdd.n62 vdd.n61 8.85536
R240 vdd.n67 vdd.n66 8.85536
R241 vdd.n352 vdd.n350 7.90638
R242 vdd.n273 vdd.n271 7.90638
R243 vdd.n194 vdd.n192 7.90638
R244 vdd.n115 vdd.n113 7.90638
R245 vdd.n41 vdd.n39 7.90638
R246 vdd.n403 vdd.n402 7.77593
R247 vdd.n458 vdd.n457 7.46309
R248 vdd.n430 vdd.n429 7.46309
R249 vdd.n461 vdd.n459 7.15344
R250 vdd.n437 vdd.n435 7.15344
R251 vdd.n412 vdd.n411 7.15344
R252 vdd.n471 vdd.n424 6.2098
R253 vdd.n447 vdd.n426 6.19834
R254 vdd.n450 vdd.n449 5.95365
R255 vdd.n420 vdd.n399 5.94964
R256 vdd.n353 vdd.t1 5.71419
R257 vdd.n274 vdd.t33 5.71419
R258 vdd.n274 vdd.t5 5.71419
R259 vdd.n195 vdd.t11 5.71419
R260 vdd.n195 vdd.t3 5.71419
R261 vdd.n116 vdd.t9 5.71419
R262 vdd.n116 vdd.t31 5.71419
R263 vdd.n42 vdd.t7 5.71419
R264 vdd.n461 vdd.n460 5.64756
R265 vdd.n437 vdd.n436 5.64756
R266 vdd.n412 vdd.n409 5.64756
R267 vdd.n149 vdd.n74 5.64054
R268 vdd.n228 vdd.n153 5.64054
R269 vdd.n307 vdd.n232 5.64054
R270 vdd.n386 vdd.n311 5.63695
R271 vdd.n71 vdd.n1 5.63695
R272 vdd.n79 vdd.n78 5.57416
R273 vdd.n158 vdd.n157 5.57416
R274 vdd.n237 vdd.n236 5.57416
R275 vdd.n432 vdd.n431 5.57212
R276 vdd.n316 vdd.n315 5.57049
R277 vdd.n405 vdd.n404 5.57042
R278 vdd.n11 vdd.n10 5.57042
R279 vdd.n388 vdd.t21 5.43072
R280 vdd.n352 vdd.n351 4.89462
R281 vdd.n273 vdd.n272 4.89462
R282 vdd.n194 vdd.n193 4.89462
R283 vdd.n115 vdd.n114 4.89462
R284 vdd.n41 vdd.n40 4.89462
R285 vdd.n388 vdd.t24 4.35663
R286 vdd.n395 vdd.t27 4.3505
R287 vdd.n395 vdd.t26 4.3505
R288 vdd.n394 vdd.t25 4.3505
R289 vdd.n394 vdd.t28 4.3505
R290 vdd.n391 vdd.t29 4.3505
R291 vdd.n391 vdd.t23 4.3505
R292 vdd.n390 vdd.t22 4.3505
R293 vdd.n390 vdd.t20 4.3505
R294 vdd.n376 vdd.n375 3.6175
R295 vdd.n370 vdd.n369 3.6175
R296 vdd.n364 vdd.n363 3.6175
R297 vdd.n358 vdd.n357 3.6175
R298 vdd.n349 vdd.n348 3.6175
R299 vdd.n344 vdd.n343 3.6175
R300 vdd.n338 vdd.n337 3.6175
R301 vdd.n332 vdd.n331 3.6175
R302 vdd.n326 vdd.n325 3.6175
R303 vdd.n320 vdd.n319 3.6175
R304 vdd.n314 vdd.n313 3.44923
R305 vdd.n297 vdd.n296 3.05241
R306 vdd.n291 vdd.n290 3.05241
R307 vdd.n285 vdd.n284 3.05241
R308 vdd.n279 vdd.n278 3.05241
R309 vdd.n270 vdd.n269 3.05241
R310 vdd.n265 vdd.n264 3.05241
R311 vdd.n259 vdd.n258 3.05241
R312 vdd.n253 vdd.n252 3.05241
R313 vdd.n247 vdd.n246 3.05241
R314 vdd.n241 vdd.n240 3.05241
R315 vdd.n218 vdd.n217 3.05241
R316 vdd.n212 vdd.n211 3.05241
R317 vdd.n206 vdd.n205 3.05241
R318 vdd.n200 vdd.n199 3.05241
R319 vdd.n191 vdd.n190 3.05241
R320 vdd.n186 vdd.n185 3.05241
R321 vdd.n180 vdd.n179 3.05241
R322 vdd.n174 vdd.n173 3.05241
R323 vdd.n168 vdd.n167 3.05241
R324 vdd.n162 vdd.n161 3.05241
R325 vdd.n139 vdd.n138 3.05241
R326 vdd.n133 vdd.n132 3.05241
R327 vdd.n127 vdd.n126 3.05241
R328 vdd.n121 vdd.n120 3.05241
R329 vdd.n112 vdd.n111 3.05241
R330 vdd.n107 vdd.n106 3.05241
R331 vdd.n101 vdd.n100 3.05241
R332 vdd.n95 vdd.n94 3.05241
R333 vdd.n89 vdd.n88 3.05241
R334 vdd.n83 vdd.n82 3.05241
R335 vdd.n235 vdd.n234 2.91084
R336 vdd.n156 vdd.n155 2.91084
R337 vdd.n77 vdd.n76 2.91084
R338 vdd.n472 vdd.n471 1.66013
R339 vdd.n150 vdd.n71 1.51623
R340 vdd.n421 vdd.n420 1.44698
R341 vdd.n450 vdd.n447 1.27483
R342 vdd.n387 vdd.n386 1.24165
R343 vdd.n308 vdd.n307 1.2194
R344 vdd.n229 vdd.n228 1.2194
R345 vdd.n150 vdd.n149 1.2194
R346 vdd.n396 vdd.n395 1.08072
R347 vdd.n392 vdd.n391 1.08072
R348 vdd.n397 vdd.n396 1.06174
R349 vdd.n393 vdd.n392 1.06174
R350 vdd.n389 vdd.n388 1.06174
R351 vdd.n433 vdd.n432 0.779301
R352 vdd.n73 vdd.n72 0.729989
R353 vdd.n152 vdd.n151 0.729989
R354 vdd.n231 vdd.n230 0.729989
R355 vdd.n407 vdd.n405 0.720048
R356 vdd.n13 vdd.n11 0.720048
R357 vdd.n318 vdd.n316 0.719967
R358 vdd.n239 vdd.n237 0.701167
R359 vdd.n160 vdd.n158 0.701167
R360 vdd.n81 vdd.n79 0.701167
R361 vdd.n423 vdd.n422 0.697387
R362 vdd.n310 vdd.n309 0.58226
R363 vdd.n7 vdd.n6 0.555728
R364 vdd.n7 vdd.n5 0.555728
R365 vdd.n7 vdd.n4 0.555728
R366 vdd.n7 vdd.n3 0.555728
R367 vdd.n7 vdd.n2 0.555728
R368 vdd.n8 vdd.n7 0.555728
R369 vdd.n421 vdd.n397 0.460436
R370 vdd.n229 vdd.n150 0.284688
R371 vdd.n308 vdd.n229 0.284688
R372 vdd.n393 vdd.n389 0.284688
R373 vdd.n397 vdd.n393 0.284688
R374 vdd.n387 vdd.n308 0.274538
R375 vdd.n472 vdd.n421 0.253438
R376 vdd vdd.n472 0.160489
R377 vdd.n447 vdd.n446 0.115891
R378 vdd.n446 vdd.n444 0.0928913
R379 vdd.n444 vdd.n441 0.0928913
R380 vdd.n441 vdd.n439 0.0928913
R381 vdd.n389 vdd.n387 0.0560556
R382 vdd.n420 vdd.n419 0.0528522
R383 vdd.n439 vdd.n438 0.0521304
R384 vdd.n386 vdd.n385 0.0519458
R385 vdd.n71 vdd.n70 0.0519458
R386 vdd.n438 vdd.n433 0.0412609
R387 vdd.n419 vdd.n417 0.0359167
R388 vdd.n417 vdd.n414 0.0359167
R389 vdd.n408 vdd.n407 0.0359167
R390 vdd.n385 vdd.n383 0.0359167
R391 vdd.n383 vdd.n380 0.0359167
R392 vdd.n380 vdd.n378 0.0359167
R393 vdd.n378 vdd.n374 0.0359167
R394 vdd.n374 vdd.n372 0.0359167
R395 vdd.n372 vdd.n368 0.0359167
R396 vdd.n368 vdd.n366 0.0359167
R397 vdd.n366 vdd.n362 0.0359167
R398 vdd.n362 vdd.n360 0.0359167
R399 vdd.n360 vdd.n356 0.0359167
R400 vdd.n356 vdd.n354 0.0359167
R401 vdd.n347 vdd.n346 0.0359167
R402 vdd.n346 vdd.n342 0.0359167
R403 vdd.n342 vdd.n340 0.0359167
R404 vdd.n340 vdd.n336 0.0359167
R405 vdd.n336 vdd.n334 0.0359167
R406 vdd.n334 vdd.n330 0.0359167
R407 vdd.n330 vdd.n328 0.0359167
R408 vdd.n328 vdd.n324 0.0359167
R409 vdd.n324 vdd.n322 0.0359167
R410 vdd.n322 vdd.n318 0.0359167
R411 vdd.n70 vdd.n68 0.0359167
R412 vdd.n68 vdd.n65 0.0359167
R413 vdd.n65 vdd.n63 0.0359167
R414 vdd.n63 vdd.n60 0.0359167
R415 vdd.n60 vdd.n58 0.0359167
R416 vdd.n58 vdd.n55 0.0359167
R417 vdd.n55 vdd.n53 0.0359167
R418 vdd.n53 vdd.n50 0.0359167
R419 vdd.n50 vdd.n48 0.0359167
R420 vdd.n48 vdd.n45 0.0359167
R421 vdd.n45 vdd.n43 0.0359167
R422 vdd.n37 vdd.n36 0.0359167
R423 vdd.n36 vdd.n33 0.0359167
R424 vdd.n33 vdd.n31 0.0359167
R425 vdd.n31 vdd.n28 0.0359167
R426 vdd.n28 vdd.n26 0.0359167
R427 vdd.n26 vdd.n23 0.0359167
R428 vdd.n23 vdd.n21 0.0359167
R429 vdd.n21 vdd.n18 0.0359167
R430 vdd.n18 vdd.n16 0.0359167
R431 vdd.n16 vdd.n13 0.0359167
R432 vdd.n452 vdd.n450 0.0330804
R433 vdd.n307 vdd.n306 0.032519
R434 vdd.n228 vdd.n227 0.032519
R435 vdd.n149 vdd.n148 0.032519
R436 vdd.n471 vdd.n470 0.0282521
R437 vdd.n470 vdd.n468 0.0224072
R438 vdd.n468 vdd.n465 0.0224072
R439 vdd.n465 vdd.n463 0.0224072
R440 vdd.n456 vdd.n455 0.0224072
R441 vdd.n455 vdd.n452 0.0224072
R442 vdd.n306 vdd.n304 0.0224072
R443 vdd.n304 vdd.n301 0.0224072
R444 vdd.n301 vdd.n299 0.0224072
R445 vdd.n299 vdd.n295 0.0224072
R446 vdd.n295 vdd.n293 0.0224072
R447 vdd.n293 vdd.n289 0.0224072
R448 vdd.n289 vdd.n287 0.0224072
R449 vdd.n287 vdd.n283 0.0224072
R450 vdd.n283 vdd.n281 0.0224072
R451 vdd.n281 vdd.n277 0.0224072
R452 vdd.n277 vdd.n275 0.0224072
R453 vdd.n268 vdd.n267 0.0224072
R454 vdd.n267 vdd.n263 0.0224072
R455 vdd.n263 vdd.n261 0.0224072
R456 vdd.n261 vdd.n257 0.0224072
R457 vdd.n257 vdd.n255 0.0224072
R458 vdd.n255 vdd.n251 0.0224072
R459 vdd.n251 vdd.n249 0.0224072
R460 vdd.n249 vdd.n245 0.0224072
R461 vdd.n245 vdd.n243 0.0224072
R462 vdd.n243 vdd.n239 0.0224072
R463 vdd.n227 vdd.n225 0.0224072
R464 vdd.n225 vdd.n222 0.0224072
R465 vdd.n222 vdd.n220 0.0224072
R466 vdd.n220 vdd.n216 0.0224072
R467 vdd.n216 vdd.n214 0.0224072
R468 vdd.n214 vdd.n210 0.0224072
R469 vdd.n210 vdd.n208 0.0224072
R470 vdd.n208 vdd.n204 0.0224072
R471 vdd.n204 vdd.n202 0.0224072
R472 vdd.n202 vdd.n198 0.0224072
R473 vdd.n198 vdd.n196 0.0224072
R474 vdd.n189 vdd.n188 0.0224072
R475 vdd.n188 vdd.n184 0.0224072
R476 vdd.n184 vdd.n182 0.0224072
R477 vdd.n182 vdd.n178 0.0224072
R478 vdd.n178 vdd.n176 0.0224072
R479 vdd.n176 vdd.n172 0.0224072
R480 vdd.n172 vdd.n170 0.0224072
R481 vdd.n170 vdd.n166 0.0224072
R482 vdd.n166 vdd.n164 0.0224072
R483 vdd.n164 vdd.n160 0.0224072
R484 vdd.n148 vdd.n146 0.0224072
R485 vdd.n146 vdd.n143 0.0224072
R486 vdd.n143 vdd.n141 0.0224072
R487 vdd.n141 vdd.n137 0.0224072
R488 vdd.n137 vdd.n135 0.0224072
R489 vdd.n135 vdd.n131 0.0224072
R490 vdd.n131 vdd.n129 0.0224072
R491 vdd.n129 vdd.n125 0.0224072
R492 vdd.n125 vdd.n123 0.0224072
R493 vdd.n123 vdd.n119 0.0224072
R494 vdd.n119 vdd.n117 0.0224072
R495 vdd.n110 vdd.n109 0.0224072
R496 vdd.n109 vdd.n105 0.0224072
R497 vdd.n105 vdd.n103 0.0224072
R498 vdd.n103 vdd.n99 0.0224072
R499 vdd.n99 vdd.n97 0.0224072
R500 vdd.n97 vdd.n93 0.0224072
R501 vdd.n93 vdd.n91 0.0224072
R502 vdd.n91 vdd.n87 0.0224072
R503 vdd.n87 vdd.n85 0.0224072
R504 vdd.n85 vdd.n81 0.0224072
R505 vdd.n354 vdd.n353 0.022375
R506 vdd.n43 vdd.n42 0.022375
R507 vdd.n413 vdd.n408 0.0202917
R508 vdd.n414 vdd.n413 0.016125
R509 vdd.n353 vdd.n347 0.0140417
R510 vdd.n42 vdd.n37 0.0140417
R511 vdd.n275 vdd.n274 0.0140309
R512 vdd.n196 vdd.n195 0.0140309
R513 vdd.n117 vdd.n116 0.0140309
R514 vdd.n463 vdd.n462 0.0127423
R515 vdd.n462 vdd.n456 0.010165
R516 vdd.n274 vdd.n268 0.00887629
R517 vdd.n195 vdd.n189 0.00887629
R518 vdd.n116 vdd.n110 0.00887629
R519 vdd.n396 vdd.n394 0.00663027
R520 vdd.n392 vdd.n390 0.00663027
R521 vdd.n438 vdd.n437 0.00190952
R522 vdd.n462 vdd.n461 0.00190952
R523 vdd.n413 vdd.n412 0.00190952
R524 vdd.n353 vdd.n352 0.00101178
R525 vdd.n274 vdd.n273 0.00101178
R526 vdd.n195 vdd.n194 0.00101178
R527 vdd.n116 vdd.n115 0.00101178
R528 vdd.n42 vdd.n41 0.00101178
R529 a_n3070_n3662.n40 a_n3070_n3662.n39 924.163
R530 a_n3070_n3662.n21 a_n3070_n3662.t13 74.7268
R531 a_n3070_n3662.n20 a_n3070_n3662.t12 74.7268
R532 a_n3070_n3662.n15 a_n3070_n3662.t14 74.7268
R533 a_n3070_n3662.n9 a_n3070_n3662.t11 74.7268
R534 a_n3070_n3662.n39 a_n3070_n3662.n0 9.3005
R535 a_n3070_n3662.n39 a_n3070_n3662.n38 9.3005
R536 a_n3070_n3662.n4 a_n3070_n3662.n1 9.10459
R537 a_n3070_n3662.n29 a_n3070_n3662.t5 4.90173
R538 a_n3070_n3662.n27 a_n3070_n3662.t9 4.90173
R539 a_n3070_n3662.n29 a_n3070_n3662.t10 4.89983
R540 a_n3070_n3662.n25 a_n3070_n3662.t1 4.89851
R541 a_n3070_n3662.n30 a_n3070_n3662.t7 4.89618
R542 a_n3070_n3662.n27 a_n3070_n3662.t4 4.89618
R543 a_n3070_n3662.n30 a_n3070_n3662.t3 4.89261
R544 a_n3070_n3662.n25 a_n3070_n3662.t6 4.89261
R545 a_n3070_n3662.n33 a_n3070_n3662.t8 4.89261
R546 a_n3070_n3662.n34 a_n3070_n3662.t2 4.36209
R547 a_n3070_n3662.n4 a_n3070_n3662.n3 3.25237
R548 a_n3070_n3662.n24 a_n3070_n3662.n18 2.7562
R549 a_n3070_n3662.n26 a_n3070_n3662.n24 1.38031
R550 a_n3070_n3662.n38 a_n3070_n3662.n37 1.30881
R551 a_n3070_n3662.n35 a_n3070_n3662.n34 1.18909
R552 a_n3070_n3662.n31 a_n3070_n3662.n30 1.07805
R553 a_n3070_n3662.n32 a_n3070_n3662.n28 1.07502
R554 a_n3070_n3662.n34 a_n3070_n3662.n33 0.538235
R555 a_n3070_n3662.n28 a_n3070_n3662.n26 0.204827
R556 a_n3070_n3662.n32 a_n3070_n3662.n31 0.204827
R557 a_n3070_n3662.n24 a_n3070_n3662.n23 0.198505
R558 a_n3070_n3662.n20 a_n3070_n3662.n19 0.16407
R559 a_n3070_n3662.n11 a_n3070_n3662.n10 0.159776
R560 a_n3070_n3662.n38 a_n3070_n3662.n4 0.0526884
R561 a_n3070_n3662.n37 a_n3070_n3662.n36 0.0426677
R562 a_n3070_n3662.n37 a_n3070_n3662.n7 0.0318735
R563 a_n3070_n3662.n17 a_n3070_n3662.n12 0.0309137
R564 a_n3070_n3662.n17 a_n3070_n3662.n16 0.0295698
R565 a_n3070_n3662.n36 a_n3070_n3662.n35 0.016125
R566 a_n3070_n3662.n22 a_n3070_n3662.n20 0.010741
R567 a_n3070_n3662.n22 a_n3070_n3662.n21 0.0107071
R568 a_n3070_n3662.n14 a_n3070_n3662.n13 0.00784719
R569 a_n3070_n3662.n7 a_n3070_n3662.n6 0.00577108
R570 a_n3070_n3662.n12 a_n3070_n3662.n11 0.00498284
R571 a_n3070_n3662.n23 a_n3070_n3662.n22 0.0040583
R572 a_n3070_n3662.n26 a_n3070_n3662.n25 0.00352842
R573 a_n3070_n3662.n28 a_n3070_n3662.n27 0.00352842
R574 a_n3070_n3662.n31 a_n3070_n3662.n29 0.00352842
R575 a_n3070_n3662.n33 a_n3070_n3662.n32 0.00352842
R576 a_n3070_n3662.n6 a_n3070_n3662.n5 0.00263488
R577 a_n3070_n3662.n9 a_n3070_n3662.n8 0.00195349
R578 a_n3070_n3662.n16 a_n3070_n3662.n15 0.00195349
R579 a_n3070_n3662.n12 a_n3070_n3662.n9 0.001503
R580 a_n3070_n3662.n3 a_n3070_n3662.n2 0.00117383
R581 a_n3070_n3662.n18 a_n3070_n3662.n17 0.00102521
R582 a_n3070_n3662.n2 a_n3070_n3662.t0 0.00101765
R583 a_n3070_n3662.n15 a_n3070_n3662.n14 0.0010022
R584 vss.n850 vss.n849 20700.8
R585 vss.t21 vss.n874 2996.99
R586 vss.n851 vss.n850 677.112
R587 vss.n877 vss.t21 634.556
R588 vss.n1000 vss.t15 449.495
R589 vss.n1000 vss.t22 449.495
R590 vss.n501 vss.t26 432.243
R591 vss.n5 vss.t5 395.844
R592 vss.n92 vss.t24 395.844
R593 vss.t7 vss.t0 310.926
R594 vss.t6 vss.t13 310.926
R595 vss.n787 vss.t28 288.082
R596 vss.n850 vss.n848 268.063
R597 vss.n316 vss.t26 245.026
R598 vss.n730 vss.t28 245.026
R599 vss.t17 vss.n315 228.767
R600 vss.n92 vss.t2 199.881
R601 vss.n93 vss.t3 199.881
R602 vss.n759 vss.n758 147.734
R603 vss.n328 vss.n327 125.654
R604 vss.n2 vss.t1 111.046
R605 vss.n8 vss.t11 100.594
R606 vss.n2 vss.t4 95.3687
R607 vss.n6 vss.t7 84.9174
R608 vss.n90 vss.t9 84.9174
R609 vss.n96 vss.t6 84.9174
R610 vss.n688 vss.n687 56.545
R611 vss.n526 vss.n524 54.4508
R612 vss.n316 vss.t17 43.9796
R613 vss.n1002 vss.t23 40.6698
R614 vss.n999 vss.t16 40.6698
R615 vss.n668 vss.t20 31.4141
R616 vss.n339 vss.n338 26.1598
R617 vss.n533 vss.n530 21.2526
R618 vss.n98 vss.n97 17.3407
R619 vss.n4 vss.n3 17.3407
R620 vss.n588 vss.n587 17.3407
R621 vss.n885 vss.n882 14.9693
R622 vss.n7 vss.n5 14.0608
R623 vss.n94 vss.n93 13.3421
R624 vss.n185 vss.n181 13.0668
R625 vss.n9 vss.n8 12.794
R626 vss.n91 vss.n90 12.794
R627 vss.n94 vss.n92 12.794
R628 vss.n7 vss.n6 12.794
R629 vss.n744 vss.t19 10.4717
R630 vss.n237 vss.n236 9.3005
R631 vss.n231 vss.n230 9.3005
R632 vss.n225 vss.n224 9.3005
R633 vss.n219 vss.n218 9.3005
R634 vss.n213 vss.n212 9.3005
R635 vss.n199 vss.n198 9.3005
R636 vss.n193 vss.n192 9.3005
R637 vss.n187 vss.n186 9.3005
R638 vss.n303 vss.n302 9.3005
R639 vss.n297 vss.n296 9.3005
R640 vss.n291 vss.n290 9.3005
R641 vss.n285 vss.n284 9.3005
R642 vss.n279 vss.n278 9.3005
R643 vss.n265 vss.n264 9.3005
R644 vss.n259 vss.n258 9.3005
R645 vss.n253 vss.n252 9.3005
R646 vss.n247 vss.n246 9.3005
R647 vss.n682 vss.n681 9.3005
R648 vss.n694 vss.n693 9.3005
R649 vss.n667 vss.n666 9.3005
R650 vss.n686 vss.n685 9.3005
R651 vss.n680 vss.n679 9.3005
R652 vss.n674 vss.n673 9.3005
R653 vss.n729 vss.n728 9.3005
R654 vss.n735 vss.n734 9.3005
R655 vss.n748 vss.n736 9.3005
R656 vss.n871 vss.n867 9.3005
R657 vss.n996 vss.n995 9.3005
R658 vss.n990 vss.n989 9.3005
R659 vss.n984 vss.n983 9.3005
R660 vss.n978 vss.n977 9.3005
R661 vss.n972 vss.n971 9.3005
R662 vss.n958 vss.n957 9.3005
R663 vss.n952 vss.n951 9.3005
R664 vss.n946 vss.n945 9.3005
R665 vss.n941 vss.n940 9.3005
R666 vss.n935 vss.n934 9.3005
R667 vss.n930 vss.n929 9.3005
R668 vss.n924 vss.n923 9.3005
R669 vss.n918 vss.n917 9.3005
R670 vss.n912 vss.n911 9.3005
R671 vss.n898 vss.n897 9.3005
R672 vss.n892 vss.n891 9.3005
R673 vss.n887 vss.n886 9.3005
R674 vss.n646 vss.n645 9.3005
R675 vss.n640 vss.n639 9.3005
R676 vss.n634 vss.n633 9.3005
R677 vss.n628 vss.n627 9.3005
R678 vss.n622 vss.n621 9.3005
R679 vss.n608 vss.n607 9.3005
R680 vss.n602 vss.n601 9.3005
R681 vss.n596 vss.n595 9.3005
R682 vss.n591 vss.n590 9.3005
R683 vss.n584 vss.n583 9.3005
R684 vss.n579 vss.n578 9.3005
R685 vss.n573 vss.n572 9.3005
R686 vss.n567 vss.n566 9.3005
R687 vss.n561 vss.n560 9.3005
R688 vss.n547 vss.n546 9.3005
R689 vss.n541 vss.n540 9.3005
R690 vss.n535 vss.n534 9.3005
R691 vss.n577 vss.n576 9.3005
R692 vss.n571 vss.n570 9.3005
R693 vss.n565 vss.n564 9.3005
R694 vss.n551 vss.n550 9.3005
R695 vss.n545 vss.n544 9.3005
R696 vss.n539 vss.n538 9.3005
R697 vss.n928 vss.n927 9.3005
R698 vss.n922 vss.n921 9.3005
R699 vss.n916 vss.n915 9.3005
R700 vss.n902 vss.n901 9.3005
R701 vss.n896 vss.n895 9.3005
R702 vss.n890 vss.n889 9.3005
R703 vss.n86 vss.n85 9.3005
R704 vss.n80 vss.n79 9.3005
R705 vss.n74 vss.n73 9.3005
R706 vss.n68 vss.n67 9.3005
R707 vss.n62 vss.n61 9.3005
R708 vss.n56 vss.n55 9.3005
R709 vss.n42 vss.n41 9.3005
R710 vss.n36 vss.n35 9.3005
R711 vss.n30 vss.n29 9.3005
R712 vss.n24 vss.n23 9.3005
R713 vss.n18 vss.n17 9.3005
R714 vss.n13 vss.n12 9.3005
R715 vss.n174 vss.n173 9.3005
R716 vss.n168 vss.n167 9.3005
R717 vss.n162 vss.n161 9.3005
R718 vss.n156 vss.n155 9.3005
R719 vss.n150 vss.n149 9.3005
R720 vss.n144 vss.n143 9.3005
R721 vss.n130 vss.n129 9.3005
R722 vss.n124 vss.n123 9.3005
R723 vss.n118 vss.n117 9.3005
R724 vss.n112 vss.n111 9.3005
R725 vss.n106 vss.n105 9.3005
R726 vss.n101 vss.n100 9.3005
R727 vss.n172 vss.n171 9.3005
R728 vss.n166 vss.n165 9.3005
R729 vss.n160 vss.n159 9.3005
R730 vss.n154 vss.n153 9.3005
R731 vss.n148 vss.n147 9.3005
R732 vss.n142 vss.n141 9.3005
R733 vss.n128 vss.n127 9.3005
R734 vss.n122 vss.n121 9.3005
R735 vss.n116 vss.n115 9.3005
R736 vss.n110 vss.n109 9.3005
R737 vss.n104 vss.n103 9.3005
R738 vss.n84 vss.n83 9.3005
R739 vss.n78 vss.n77 9.3005
R740 vss.n72 vss.n71 9.3005
R741 vss.n66 vss.n65 9.3005
R742 vss.n60 vss.n59 9.3005
R743 vss.n54 vss.n53 9.3005
R744 vss.n40 vss.n39 9.3005
R745 vss.n34 vss.n33 9.3005
R746 vss.n28 vss.n27 9.3005
R747 vss.n22 vss.n21 9.3005
R748 vss.n16 vss.n15 9.3005
R749 vss.n301 vss.n300 9.3005
R750 vss.n295 vss.n294 9.3005
R751 vss.n289 vss.n288 9.3005
R752 vss.n283 vss.n282 9.3005
R753 vss.n269 vss.n268 9.3005
R754 vss.n263 vss.n262 9.3005
R755 vss.n257 vss.n256 9.3005
R756 vss.n251 vss.n250 9.3005
R757 vss.n235 vss.n234 9.3005
R758 vss.n229 vss.n228 9.3005
R759 vss.n223 vss.n222 9.3005
R760 vss.n217 vss.n216 9.3005
R761 vss.n203 vss.n202 9.3005
R762 vss.n197 vss.n196 9.3005
R763 vss.n191 vss.n190 9.3005
R764 vss.n321 vss.n320 9.3005
R765 vss.n314 vss.n313 9.3005
R766 vss.n384 vss.n383 9.3005
R767 vss.n390 vss.n389 9.3005
R768 vss.n336 vss.n335 9.3005
R769 vss.n403 vss.n391 9.3005
R770 vss.n521 vss.n489 9.3005
R771 vss.n994 vss.n993 9.3005
R772 vss.n988 vss.n987 9.3005
R773 vss.n982 vss.n981 9.3005
R774 vss.n976 vss.n975 9.3005
R775 vss.n962 vss.n961 9.3005
R776 vss.n956 vss.n955 9.3005
R777 vss.n950 vss.n949 9.3005
R778 vss.n944 vss.n943 9.3005
R779 vss.n388 vss.n387 9.3005
R780 vss.n319 vss.n318 9.3005
R781 vss.n644 vss.n643 9.3005
R782 vss.n638 vss.n637 9.3005
R783 vss.n632 vss.n631 9.3005
R784 vss.n626 vss.n625 9.3005
R785 vss.n612 vss.n611 9.3005
R786 vss.n606 vss.n605 9.3005
R787 vss.n600 vss.n599 9.3005
R788 vss.n594 vss.n593 9.3005
R789 vss.n582 vss.n581 9.3005
R790 vss.n733 vss.n732 9.3005
R791 vss.n678 vss.n677 9.3005
R792 vss.n691 vss.n690 9.3005
R793 vss.n671 vss.n670 9.3005
R794 vss.n933 vss.n932 9.3005
R795 vss.n832 vss.n831 9.15497
R796 vss.n831 vss.n830 9.15497
R797 vss.n761 vss.n760 9.15497
R798 vss.n760 vss.n759 9.15497
R799 vss.n773 vss.n772 9.15497
R800 vss.n772 vss.n771 9.15497
R801 vss.n789 vss.n788 9.15497
R802 vss.n788 vss.n787 9.15497
R803 vss.n816 vss.n815 9.15497
R804 vss.n815 vss.n814 9.15497
R805 vss.n854 vss.n853 9.15497
R806 vss.n857 vss.n856 9.15497
R807 vss.n829 vss.n828 9.15497
R808 vss.n846 vss.n845 9.15497
R809 vss.n845 vss.n844 9.15497
R810 vss.n861 vss.n860 9.15497
R811 vss.n860 vss.n859 9.15497
R812 vss.n842 vss.n841 9.15497
R813 vss.n841 vss.n840 9.15497
R814 vss.n865 vss.n864 9.15497
R815 vss.n864 vss.n863 9.15497
R816 vss.n838 vss.n837 9.15497
R817 vss.n837 vss.n836 9.15497
R818 vss.n870 vss.n869 9.15497
R819 vss.n576 vss.n575 9.15497
R820 vss.n570 vss.n569 9.15497
R821 vss.n564 vss.n563 9.15497
R822 vss.n556 vss.n555 9.15497
R823 vss.n550 vss.n549 9.15497
R824 vss.n544 vss.n543 9.15497
R825 vss.n538 vss.n537 9.15497
R826 vss.n532 vss.n531 9.15497
R827 vss.n927 vss.n926 9.15497
R828 vss.n921 vss.n920 9.15497
R829 vss.n915 vss.n914 9.15497
R830 vss.n907 vss.n906 9.15497
R831 vss.n901 vss.n900 9.15497
R832 vss.n895 vss.n894 9.15497
R833 vss.n889 vss.n888 9.15497
R834 vss.n884 vss.n883 9.15497
R835 vss.n171 vss.n170 9.15497
R836 vss.n165 vss.n164 9.15497
R837 vss.n159 vss.n158 9.15497
R838 vss.n153 vss.n152 9.15497
R839 vss.n147 vss.n146 9.15497
R840 vss.n141 vss.n140 9.15497
R841 vss.n134 vss.n133 9.15497
R842 vss.n127 vss.n126 9.15497
R843 vss.n121 vss.n120 9.15497
R844 vss.n115 vss.n114 9.15497
R845 vss.n109 vss.n108 9.15497
R846 vss.n103 vss.n102 9.15497
R847 vss.n89 vss.n88 9.15497
R848 vss.n83 vss.n82 9.15497
R849 vss.n77 vss.n76 9.15497
R850 vss.n71 vss.n70 9.15497
R851 vss.n65 vss.n64 9.15497
R852 vss.n59 vss.n58 9.15497
R853 vss.n53 vss.n52 9.15497
R854 vss.n46 vss.n45 9.15497
R855 vss.n39 vss.n38 9.15497
R856 vss.n33 vss.n32 9.15497
R857 vss.n27 vss.n26 9.15497
R858 vss.n21 vss.n20 9.15497
R859 vss.n15 vss.n14 9.15497
R860 vss.n1 vss.n0 9.15497
R861 vss.n300 vss.n299 9.15497
R862 vss.n299 vss.n298 9.15497
R863 vss.n294 vss.n293 9.15497
R864 vss.n293 vss.n292 9.15497
R865 vss.n288 vss.n287 9.15497
R866 vss.n287 vss.n286 9.15497
R867 vss.n282 vss.n281 9.15497
R868 vss.n281 vss.n280 9.15497
R869 vss.n274 vss.n273 9.15497
R870 vss.n273 vss.n272 9.15497
R871 vss.n268 vss.n267 9.15497
R872 vss.n267 vss.n266 9.15497
R873 vss.n262 vss.n261 9.15497
R874 vss.n261 vss.n260 9.15497
R875 vss.n256 vss.n255 9.15497
R876 vss.n255 vss.n254 9.15497
R877 vss.n250 vss.n249 9.15497
R878 vss.n249 vss.n248 9.15497
R879 vss.n244 vss.n243 9.15497
R880 vss.n243 vss.n242 9.15497
R881 vss.n179 vss.n178 9.15497
R882 vss.n178 vss.n177 9.15497
R883 vss.n234 vss.n233 9.15497
R884 vss.n233 vss.n232 9.15497
R885 vss.n228 vss.n227 9.15497
R886 vss.n227 vss.n226 9.15497
R887 vss.n222 vss.n221 9.15497
R888 vss.n221 vss.n220 9.15497
R889 vss.n216 vss.n215 9.15497
R890 vss.n215 vss.n214 9.15497
R891 vss.n208 vss.n207 9.15497
R892 vss.n207 vss.n206 9.15497
R893 vss.n202 vss.n201 9.15497
R894 vss.n201 vss.n200 9.15497
R895 vss.n196 vss.n195 9.15497
R896 vss.n195 vss.n194 9.15497
R897 vss.n190 vss.n189 9.15497
R898 vss.n189 vss.n188 9.15497
R899 vss.n184 vss.n183 9.15497
R900 vss.n183 vss.n182 9.15497
R901 vss.n181 vss.n180 9.15497
R902 vss.n240 vss.n239 9.15497
R903 vss.n239 vss.n238 9.15497
R904 vss.n341 vss.n340 9.15497
R905 vss.n340 vss.n339 9.15497
R906 vss.n333 vss.n332 9.15497
R907 vss.n348 vss.n347 9.15497
R908 vss.n347 vss.n346 9.15497
R909 vss.n361 vss.n360 9.15497
R910 vss.n360 vss.n359 9.15497
R911 vss.n379 vss.n378 9.15497
R912 vss.n378 vss.n377 9.15497
R913 vss.n326 vss.n325 9.15497
R914 vss.n481 vss.n480 9.15497
R915 vss.n480 vss.n479 9.15497
R916 vss.n469 vss.n468 9.15497
R917 vss.n468 vss.n467 9.15497
R918 vss.n514 vss.n513 9.15497
R919 vss.n511 vss.n510 9.15497
R920 vss.n510 vss.n509 9.15497
R921 vss.n507 vss.n506 9.15497
R922 vss.n506 vss.n505 9.15497
R923 vss.n503 vss.n502 9.15497
R924 vss.n502 vss.n501 9.15497
R925 vss.n499 vss.n498 9.15497
R926 vss.n498 vss.n497 9.15497
R927 vss.n495 vss.n494 9.15497
R928 vss.n494 vss.n493 9.15497
R929 vss.n491 vss.n490 9.15497
R930 vss.n520 vss.n519 9.15497
R931 vss.n485 vss.n484 9.15497
R932 vss.n473 vss.n472 9.15497
R933 vss.n414 vss.n413 9.15497
R934 vss.n426 vss.n425 9.15497
R935 vss.n441 vss.n440 9.15497
R936 vss.n661 vss.n660 9.15497
R937 vss.n699 vss.n698 9.15497
R938 vss.n719 vss.n718 9.15497
R939 vss.n820 vss.n819 9.15497
R940 vss.n993 vss.n992 9.15497
R941 vss.n987 vss.n986 9.15497
R942 vss.n981 vss.n980 9.15497
R943 vss.n975 vss.n974 9.15497
R944 vss.n967 vss.n966 9.15497
R945 vss.n961 vss.n960 9.15497
R946 vss.n955 vss.n954 9.15497
R947 vss.n949 vss.n948 9.15497
R948 vss.n943 vss.n942 9.15497
R949 vss.n879 vss.n878 9.15497
R950 vss.n878 vss.n877 9.15497
R951 vss.n330 vss.n329 9.15497
R952 vss.n329 vss.n328 9.15497
R953 vss.n318 vss.n317 9.15497
R954 vss.n317 vss.n316 9.15497
R955 vss.n387 vss.n386 9.15497
R956 vss.n386 vss.n385 9.15497
R957 vss.n394 vss.n393 9.15497
R958 vss.n393 vss.n392 9.15497
R959 vss.n401 vss.n400 9.15497
R960 vss.n400 vss.n399 9.15497
R961 vss.n398 vss.n397 9.15497
R962 vss.n408 vss.n407 9.15497
R963 vss.n643 vss.n642 9.15497
R964 vss.n637 vss.n636 9.15497
R965 vss.n631 vss.n630 9.15497
R966 vss.n625 vss.n624 9.15497
R967 vss.n617 vss.n616 9.15497
R968 vss.n611 vss.n610 9.15497
R969 vss.n605 vss.n604 9.15497
R970 vss.n599 vss.n598 9.15497
R971 vss.n593 vss.n592 9.15497
R972 vss.n528 vss.n527 9.15497
R973 vss.n527 vss.n526 9.15497
R974 vss.n581 vss.n580 9.15497
R975 vss.n670 vss.n669 9.15497
R976 vss.n669 vss.n668 9.15497
R977 vss.n690 vss.n689 9.15497
R978 vss.n689 vss.n688 9.15497
R979 vss.n677 vss.n676 9.15497
R980 vss.n676 vss.n675 9.15497
R981 vss.n732 vss.n731 9.15497
R982 vss.n731 vss.n730 9.15497
R983 vss.n746 vss.n745 9.15497
R984 vss.n745 vss.n744 9.15497
R985 vss.n739 vss.n738 9.15497
R986 vss.n738 vss.n737 9.15497
R987 vss.n742 vss.n741 9.15497
R988 vss.n659 vss.n658 9.15497
R989 vss.n753 vss.n752 9.15497
R990 vss.n655 vss.n654 9.15497
R991 vss.n932 vss.n931 9.15497
R992 vss.n438 vss.n437 8.85536
R993 vss.n785 vss.n784 8.85536
R994 vss.n685 vss.n684 8.85536
R995 vss.n673 vss.n672 8.85536
R996 vss.n728 vss.n727 8.85536
R997 vss.n716 vss.n715 8.85536
R998 vss.n704 vss.n703 8.85536
R999 vss.n764 vss.n763 8.85536
R1000 vss.n776 vss.n775 8.85536
R1001 vss.n801 vss.n800 8.85536
R1002 vss.n798 vss.n797 8.85536
R1003 vss.n805 vss.n804 8.85536
R1004 vss.n808 vss.n807 8.85536
R1005 vss.n313 vss.n312 8.85536
R1006 vss.n383 vss.n382 8.85536
R1007 vss.n352 vss.n351 8.85536
R1008 vss.n375 vss.n374 8.85536
R1009 vss.n364 vss.n363 8.85536
R1010 vss.n417 vss.n416 8.85536
R1011 vss.n429 vss.n428 8.85536
R1012 vss.n453 vss.n452 8.85536
R1013 vss.n450 vss.n449 8.85536
R1014 vss.n457 vss.n456 8.85536
R1015 vss.n461 vss.n460 8.85536
R1016 vss.n784 vss.n783 8.40958
R1017 vss.n437 vss.n436 8.40958
R1018 vss.n374 vss.n373 8.3985
R1019 vss.n715 vss.n714 8.3985
R1020 vss.n853 vss.n852 8.04597
R1021 vss.n519 vss.n518 8.04553
R1022 vss.n698 vss.n697 8.04553
R1023 vss.n819 vss.n818 8.04553
R1024 vss.n325 vss.n324 8.04506
R1025 vss.n472 vss.n471 8.04503
R1026 vss.n425 vss.n424 8.04503
R1027 vss.n48 vss.n46 7.90638
R1028 vss.n136 vss.n134 7.90638
R1029 vss.n209 vss.n205 7.15344
R1030 vss.n275 vss.n271 7.15344
R1031 vss.n968 vss.n964 7.15344
R1032 vss.n908 vss.n904 7.15344
R1033 vss.n618 vss.n614 7.15344
R1034 vss.n557 vss.n553 7.15344
R1035 vss.n882 vss.n881 7.14271
R1036 vss.n460 vss.n459 7.0309
R1037 vss.n1001 vss.n1000 6.88684
R1038 vss.n175 vss.n89 6.2098
R1039 vss.n87 vss.n1 6.2098
R1040 vss.n304 vss.n179 6.19834
R1041 vss.n997 vss.n879 6.19834
R1042 vss.n647 vss.n528 6.19834
R1043 vss.n241 vss.n240 6.19834
R1044 vss.n937 vss.n936 6.19834
R1045 vss.n586 vss.n585 6.19834
R1046 vss.n484 vss.n483 6.1288
R1047 vss.n407 vss.n406 6.1288
R1048 vss.n752 vss.n751 6.1288
R1049 vss.n658 vss.n657 6.01858
R1050 vss.n828 vss.n827 6.01829
R1051 vss.n245 vss.n244 5.73064
R1052 vss.n939 vss.n938 5.73064
R1053 vss.n589 vss.n588 5.73064
R1054 vss.n843 vss.n842 5.71564
R1055 vss.n500 vss.n499 5.71564
R1056 vss.n209 vss.n208 5.64756
R1057 vss.n275 vss.n274 5.64756
R1058 vss.n968 vss.n967 5.64756
R1059 vss.n908 vss.n907 5.64756
R1060 vss.n618 vss.n617 5.64756
R1061 vss.n557 vss.n556 5.64756
R1062 vss.n11 vss.n4 5.64054
R1063 vss.n99 vss.n98 5.64054
R1064 vss.n185 vss.n184 5.58665
R1065 vss.n885 vss.n884 5.58665
R1066 vss.n533 vss.n532 5.58665
R1067 vss.n871 vss.n870 5.28049
R1068 vss.n336 vss.n326 5.28049
R1069 vss.n521 vss.n520 5.28049
R1070 vss.n464 vss.n455 5.25157
R1071 vss.n420 vss.n419 5.25157
R1072 vss.n811 vss.n803 5.25157
R1073 vss.n767 vss.n766 5.25157
R1074 vss.n871 vss.n855 5.25007
R1075 vss.n748 vss.n743 5.25007
R1076 vss.n521 vss.n515 5.25007
R1077 vss.n811 vss.n810 5.22057
R1078 vss.n355 vss.n354 5.22057
R1079 vss.n464 vss.n463 5.20217
R1080 vss.n704 vss.n702 5.15606
R1081 vss.n305 vss.n304 5.12896
R1082 vss.n998 vss.n997 5.12896
R1083 vss.n648 vss.n647 5.12896
R1084 vss.n48 vss.n47 4.89462
R1085 vss.n136 vss.n135 4.89462
R1086 vss.n662 vss.n659 4.30941
R1087 vss.n662 vss.n661 4.30941
R1088 vss.n748 vss.n740 3.77639
R1089 vss.n748 vss.n747 3.77639
R1090 vss.n871 vss.n858 3.77639
R1091 vss.n871 vss.n847 3.77639
R1092 vss.n871 vss.n862 3.77639
R1093 vss.n871 vss.n866 3.77639
R1094 vss.n871 vss.n839 3.77639
R1095 vss.n336 vss.n331 3.77639
R1096 vss.n336 vss.n334 3.77639
R1097 vss.n403 vss.n395 3.77639
R1098 vss.n521 vss.n512 3.77639
R1099 vss.n521 vss.n508 3.77639
R1100 vss.n521 vss.n504 3.77639
R1101 vss.n521 vss.n496 3.77639
R1102 vss.n521 vss.n492 3.77639
R1103 vss.n811 vss.n799 3.51051
R1104 vss.n811 vss.n806 3.51051
R1105 vss.n464 vss.n451 3.51051
R1106 vss.n464 vss.n458 3.51051
R1107 vss.n137 vss.t14 3.48118
R1108 vss.n137 vss.t10 3.48118
R1109 vss.n49 vss.t8 3.48118
R1110 vss.n49 vss.t12 3.48118
R1111 vss.n717 vss.n716 3.1005
R1112 vss.n705 vss.n704 3.1005
R1113 vss.n786 vss.n785 3.1005
R1114 vss.n777 vss.n776 3.1005
R1115 vss.n833 vss.n829 3.1005
R1116 vss.n833 vss.n832 3.1005
R1117 vss.n762 vss.n761 3.1005
R1118 vss.n774 vss.n773 3.1005
R1119 vss.n790 vss.n789 3.1005
R1120 vss.n821 vss.n816 3.1005
R1121 vss.n342 vss.n341 3.1005
R1122 vss.n349 vss.n348 3.1005
R1123 vss.n362 vss.n361 3.1005
R1124 vss.n380 vss.n379 3.1005
R1125 vss.n376 vss.n375 3.1005
R1126 vss.n365 vss.n364 3.1005
R1127 vss.n439 vss.n438 3.1005
R1128 vss.n430 vss.n429 3.1005
R1129 vss.n486 vss.n481 3.1005
R1130 vss.n474 vss.n469 3.1005
R1131 vss.n486 vss.n485 3.1005
R1132 vss.n474 vss.n473 3.1005
R1133 vss.n415 vss.n414 3.1005
R1134 vss.n427 vss.n426 3.1005
R1135 vss.n442 vss.n441 3.1005
R1136 vss.n700 vss.n699 3.1005
R1137 vss.n720 vss.n719 3.1005
R1138 vss.n821 vss.n820 3.1005
R1139 vss.n409 vss.n408 3.1005
R1140 vss.n754 vss.n753 3.1005
R1141 vss.n402 vss.n401 2.9463
R1142 vss.n402 vss.n398 2.94569
R1143 vss.n948 vss.n947 2.42332
R1144 vss.n954 vss.n953 2.42332
R1145 vss.n960 vss.n959 2.42332
R1146 vss.n966 vss.n965 2.42332
R1147 vss.n974 vss.n973 2.42332
R1148 vss.n980 vss.n979 2.42332
R1149 vss.n986 vss.n985 2.42332
R1150 vss.n992 vss.n991 2.38585
R1151 vss.n351 vss.n350 2.35017
R1152 vss.n684 vss.n683 2.35017
R1153 vss.n245 vss.n241 2.31211
R1154 vss.n939 vss.n937 2.31211
R1155 vss.n589 vss.n586 2.31211
R1156 vss.n458 vss.n457 2.28197
R1157 vss.n806 vss.n805 2.28197
R1158 vss.n799 vss.n798 2.28197
R1159 vss.n451 vss.n450 2.28197
R1160 vss.n659 vss.n655 2.28169
R1161 vss.n405 vss.t18 2.09474
R1162 vss.n598 vss.n597 1.93234
R1163 vss.n604 vss.n603 1.93234
R1164 vss.n610 vss.n609 1.93234
R1165 vss.n616 vss.n615 1.93234
R1166 vss.n624 vss.n623 1.93234
R1167 vss.n630 vss.n629 1.93234
R1168 vss.n636 vss.n635 1.93234
R1169 vss.n894 vss.n893 1.93234
R1170 vss.n900 vss.n899 1.93234
R1171 vss.n906 vss.n905 1.93234
R1172 vss.n914 vss.n913 1.93234
R1173 vss.n920 vss.n919 1.93234
R1174 vss.n537 vss.n536 1.93234
R1175 vss.n543 vss.n542 1.93234
R1176 vss.n549 vss.n548 1.93234
R1177 vss.n555 vss.n554 1.93234
R1178 vss.n563 vss.n562 1.93234
R1179 vss.n569 vss.n568 1.93234
R1180 vss.n20 vss.n19 1.93234
R1181 vss.n26 vss.n25 1.93234
R1182 vss.n32 vss.n31 1.93234
R1183 vss.n38 vss.n37 1.93234
R1184 vss.n45 vss.n44 1.93234
R1185 vss.n52 vss.n51 1.93234
R1186 vss.n58 vss.n57 1.93234
R1187 vss.n64 vss.n63 1.93234
R1188 vss.n70 vss.n69 1.93234
R1189 vss.n76 vss.n75 1.93234
R1190 vss.n108 vss.n107 1.93234
R1191 vss.n114 vss.n113 1.93234
R1192 vss.n120 vss.n119 1.93234
R1193 vss.n126 vss.n125 1.93234
R1194 vss.n133 vss.n132 1.93234
R1195 vss.n140 vss.n139 1.93234
R1196 vss.n146 vss.n145 1.93234
R1197 vss.n152 vss.n151 1.93234
R1198 vss.n158 vss.n157 1.93234
R1199 vss.n164 vss.n163 1.93234
R1200 vss.n419 vss.n418 1.92507
R1201 vss.n766 vss.n765 1.92507
R1202 vss.n354 vss.n353 1.92211
R1203 vss.n642 vss.n641 1.90249
R1204 vss.n926 vss.n925 1.90249
R1205 vss.n575 vss.n574 1.90249
R1206 vss.n82 vss.n81 1.90249
R1207 vss.n170 vss.n169 1.90249
R1208 vss.n403 vss.n402 1.8362
R1209 vss.n858 vss.n857 1.75023
R1210 vss.n847 vss.n846 1.75023
R1211 vss.n862 vss.n861 1.75023
R1212 vss.n866 vss.n865 1.75023
R1213 vss.n839 vss.n838 1.75023
R1214 vss.n334 vss.n333 1.75023
R1215 vss.n512 vss.n511 1.75023
R1216 vss.n508 vss.n507 1.75023
R1217 vss.n504 vss.n503 1.75023
R1218 vss.n496 vss.n495 1.75023
R1219 vss.n492 vss.n491 1.75023
R1220 vss.n395 vss.n394 1.75023
R1221 vss.n331 vss.n330 1.75023
R1222 vss.n740 vss.n739 1.75023
R1223 vss.n747 vss.n746 1.75023
R1224 vss.n827 vss.n826 1.57034
R1225 vss.n657 vss.n656 1.56991
R1226 vss.n483 vss.n482 1.51507
R1227 vss.n406 vss.n405 1.51507
R1228 vss.n751 vss.n750 1.51507
R1229 vss.n702 vss.n701 1.42272
R1230 vss.n455 vss.n454 1.21396
R1231 vss.n803 vss.n802 1.21396
R1232 vss.n810 vss.n809 1.21099
R1233 vss.n176 vss.n87 0.995287
R1234 vss.n95 vss.n94 0.993288
R1235 vss.n187 vss.n185 0.762358
R1236 vss.n887 vss.n885 0.762358
R1237 vss.n535 vss.n533 0.762358
R1238 vss.n176 vss.n175 0.711099
R1239 vss.n463 vss.n462 0.656018
R1240 vss.n305 vss.n176 0.612145
R1241 vss.n11 vss.n10 0.607836
R1242 vss.n99 vss.n95 0.607836
R1243 vss.t27 vss.n711 0.599391
R1244 vss.t27 vss.n712 0.599391
R1245 vss.t25 vss.n371 0.599391
R1246 vss.t25 vss.n372 0.599391
R1247 vss.t27 vss.n713 0.599342
R1248 vss.n518 vss.n517 0.556698
R1249 vss.n818 vss.n817 0.556698
R1250 vss.n852 vss.n851 0.556239
R1251 vss.n471 vss.n470 0.556239
R1252 vss.n324 vss.n323 0.556206
R1253 vss.n881 vss.n880 0.497022
R1254 vss.n530 vss.n529 0.490159
R1255 vss.n97 vss.n96 0.490159
R1256 vss.n3 vss.n2 0.490159
R1257 vss.n526 vss.n525 0.482453
R1258 vss.n877 vss.n876 0.482453
R1259 vss.n999 vss.n998 0.430788
R1260 vss.n877 vss.n875 0.37528
R1261 vss.n354 vss.n352 0.356981
R1262 vss.n810 vss.n808 0.356981
R1263 vss.n766 vss.n764 0.354276
R1264 vss.n803 vss.n801 0.354276
R1265 vss.n419 vss.n417 0.354276
R1266 vss.n455 vss.n453 0.354276
R1267 vss.n463 vss.n461 0.345484
R1268 vss.n10 vss.n7 0.286558
R1269 vss.n95 vss.n91 0.286558
R1270 vss.n10 vss.n9 0.272135
R1271 vss.n870 vss.n868 0.253965
R1272 vss.n655 vss.n653 0.253965
R1273 vss.n326 vss.n322 0.253965
R1274 vss.n520 vss.n516 0.253965
R1275 vss.n714 vss.t27 0.23529
R1276 vss.n373 vss.t25 0.23529
R1277 vss.n648 vss.n523 0.165831
R1278 vss.n873 vss.n648 0.154079
R1279 vss.n873 vss.n872 0.151997
R1280 vss.n523 vss.n522 0.151997
R1281 vss.n1002 vss.n1001 0.143662
R1282 vss.n1001 vss.n999 0.141526
R1283 vss.n247 vss.n245 0.134638
R1284 vss.n941 vss.n939 0.134638
R1285 vss.n591 vss.n589 0.134638
R1286 vss.n998 vss.n873 0.131109
R1287 vss.n398 vss.n396 0.127233
R1288 vss.n523 vss.n305 0.119357
R1289 vss.n241 vss.n237 0.115891
R1290 vss.n304 vss.n303 0.115891
R1291 vss.n937 vss.n935 0.115891
R1292 vss.n997 vss.n996 0.115891
R1293 vss.n586 vss.n584 0.115891
R1294 vss.n647 vss.n646 0.115891
R1295 vss.n191 vss.n187 0.0928913
R1296 vss.n193 vss.n191 0.0928913
R1297 vss.n197 vss.n193 0.0928913
R1298 vss.n199 vss.n197 0.0928913
R1299 vss.n203 vss.n199 0.0928913
R1300 vss.n204 vss.n203 0.0928913
R1301 vss.n213 vss.n211 0.0928913
R1302 vss.n217 vss.n213 0.0928913
R1303 vss.n219 vss.n217 0.0928913
R1304 vss.n223 vss.n219 0.0928913
R1305 vss.n225 vss.n223 0.0928913
R1306 vss.n229 vss.n225 0.0928913
R1307 vss.n231 vss.n229 0.0928913
R1308 vss.n235 vss.n231 0.0928913
R1309 vss.n237 vss.n235 0.0928913
R1310 vss.n251 vss.n247 0.0928913
R1311 vss.n253 vss.n251 0.0928913
R1312 vss.n257 vss.n253 0.0928913
R1313 vss.n259 vss.n257 0.0928913
R1314 vss.n263 vss.n259 0.0928913
R1315 vss.n265 vss.n263 0.0928913
R1316 vss.n269 vss.n265 0.0928913
R1317 vss.n270 vss.n269 0.0928913
R1318 vss.n279 vss.n277 0.0928913
R1319 vss.n283 vss.n279 0.0928913
R1320 vss.n285 vss.n283 0.0928913
R1321 vss.n289 vss.n285 0.0928913
R1322 vss.n291 vss.n289 0.0928913
R1323 vss.n295 vss.n291 0.0928913
R1324 vss.n297 vss.n295 0.0928913
R1325 vss.n301 vss.n297 0.0928913
R1326 vss.n303 vss.n301 0.0928913
R1327 vss.n890 vss.n887 0.0928913
R1328 vss.n892 vss.n890 0.0928913
R1329 vss.n896 vss.n892 0.0928913
R1330 vss.n898 vss.n896 0.0928913
R1331 vss.n902 vss.n898 0.0928913
R1332 vss.n903 vss.n902 0.0928913
R1333 vss.n912 vss.n910 0.0928913
R1334 vss.n916 vss.n912 0.0928913
R1335 vss.n918 vss.n916 0.0928913
R1336 vss.n922 vss.n918 0.0928913
R1337 vss.n924 vss.n922 0.0928913
R1338 vss.n928 vss.n924 0.0928913
R1339 vss.n930 vss.n928 0.0928913
R1340 vss.n933 vss.n930 0.0928913
R1341 vss.n935 vss.n933 0.0928913
R1342 vss.n944 vss.n941 0.0928913
R1343 vss.n946 vss.n944 0.0928913
R1344 vss.n950 vss.n946 0.0928913
R1345 vss.n952 vss.n950 0.0928913
R1346 vss.n956 vss.n952 0.0928913
R1347 vss.n958 vss.n956 0.0928913
R1348 vss.n962 vss.n958 0.0928913
R1349 vss.n963 vss.n962 0.0928913
R1350 vss.n972 vss.n970 0.0928913
R1351 vss.n976 vss.n972 0.0928913
R1352 vss.n978 vss.n976 0.0928913
R1353 vss.n982 vss.n978 0.0928913
R1354 vss.n984 vss.n982 0.0928913
R1355 vss.n988 vss.n984 0.0928913
R1356 vss.n990 vss.n988 0.0928913
R1357 vss.n994 vss.n990 0.0928913
R1358 vss.n996 vss.n994 0.0928913
R1359 vss.n539 vss.n535 0.0928913
R1360 vss.n541 vss.n539 0.0928913
R1361 vss.n545 vss.n541 0.0928913
R1362 vss.n547 vss.n545 0.0928913
R1363 vss.n551 vss.n547 0.0928913
R1364 vss.n552 vss.n551 0.0928913
R1365 vss.n561 vss.n559 0.0928913
R1366 vss.n565 vss.n561 0.0928913
R1367 vss.n567 vss.n565 0.0928913
R1368 vss.n571 vss.n567 0.0928913
R1369 vss.n573 vss.n571 0.0928913
R1370 vss.n577 vss.n573 0.0928913
R1371 vss.n579 vss.n577 0.0928913
R1372 vss.n582 vss.n579 0.0928913
R1373 vss.n584 vss.n582 0.0928913
R1374 vss.n594 vss.n591 0.0928913
R1375 vss.n596 vss.n594 0.0928913
R1376 vss.n600 vss.n596 0.0928913
R1377 vss.n602 vss.n600 0.0928913
R1378 vss.n606 vss.n602 0.0928913
R1379 vss.n608 vss.n606 0.0928913
R1380 vss.n612 vss.n608 0.0928913
R1381 vss.n613 vss.n612 0.0928913
R1382 vss.n622 vss.n620 0.0928913
R1383 vss.n626 vss.n622 0.0928913
R1384 vss.n628 vss.n626 0.0928913
R1385 vss.n632 vss.n628 0.0928913
R1386 vss.n634 vss.n632 0.0928913
R1387 vss.n638 vss.n634 0.0928913
R1388 vss.n640 vss.n638 0.0928913
R1389 vss.n644 vss.n640 0.0928913
R1390 vss.n646 vss.n644 0.0928913
R1391 vss.n708 vss.n705 0.0568063
R1392 vss.n314 vss.n311 0.0568063
R1393 vss.n780 vss.n777 0.0563036
R1394 vss.n433 vss.n430 0.0563036
R1395 vss.n729 vss.n726 0.0562432
R1396 vss.n368 vss.n365 0.0558097
R1397 vss.n855 vss.n854 0.0554606
R1398 vss.n515 vss.n514 0.0554606
R1399 vss.n743 vss.n742 0.0554606
R1400 vss.n717 vss.n710 0.0551171
R1401 vss.n786 vss.n782 0.0546295
R1402 vss.n439 vss.n435 0.0546295
R1403 vss.n376 vss.n370 0.0541504
R1404 vss.n210 vss.n204 0.0521304
R1405 vss.n276 vss.n270 0.0521304
R1406 vss.n909 vss.n903 0.0521304
R1407 vss.n969 vss.n963 0.0521304
R1408 vss.n558 vss.n552 0.0521304
R1409 vss.n619 vss.n613 0.0521304
R1410 vss.n211 vss.n210 0.0412609
R1411 vss.n277 vss.n276 0.0412609
R1412 vss.n910 vss.n909 0.0412609
R1413 vss.n970 vss.n969 0.0412609
R1414 vss.n559 vss.n558 0.0412609
R1415 vss.n620 vss.n619 0.0412609
R1416 vss.n13 vss.n11 0.032519
R1417 vss.n101 vss.n99 0.032519
R1418 vss.n87 vss.n86 0.0282521
R1419 vss.n175 vss.n174 0.0282521
R1420 vss.n749 vss.n748 0.0228214
R1421 vss.n404 vss.n403 0.0228214
R1422 vss.n337 vss.n336 0.0226239
R1423 vss.n16 vss.n13 0.0224072
R1424 vss.n18 vss.n16 0.0224072
R1425 vss.n22 vss.n18 0.0224072
R1426 vss.n24 vss.n22 0.0224072
R1427 vss.n28 vss.n24 0.0224072
R1428 vss.n30 vss.n28 0.0224072
R1429 vss.n34 vss.n30 0.0224072
R1430 vss.n36 vss.n34 0.0224072
R1431 vss.n40 vss.n36 0.0224072
R1432 vss.n42 vss.n40 0.0224072
R1433 vss.n43 vss.n42 0.0224072
R1434 vss.n54 vss.n50 0.0224072
R1435 vss.n56 vss.n54 0.0224072
R1436 vss.n60 vss.n56 0.0224072
R1437 vss.n62 vss.n60 0.0224072
R1438 vss.n66 vss.n62 0.0224072
R1439 vss.n68 vss.n66 0.0224072
R1440 vss.n72 vss.n68 0.0224072
R1441 vss.n74 vss.n72 0.0224072
R1442 vss.n78 vss.n74 0.0224072
R1443 vss.n80 vss.n78 0.0224072
R1444 vss.n84 vss.n80 0.0224072
R1445 vss.n86 vss.n84 0.0224072
R1446 vss.n104 vss.n101 0.0224072
R1447 vss.n106 vss.n104 0.0224072
R1448 vss.n110 vss.n106 0.0224072
R1449 vss.n112 vss.n110 0.0224072
R1450 vss.n116 vss.n112 0.0224072
R1451 vss.n118 vss.n116 0.0224072
R1452 vss.n122 vss.n118 0.0224072
R1453 vss.n124 vss.n122 0.0224072
R1454 vss.n128 vss.n124 0.0224072
R1455 vss.n130 vss.n128 0.0224072
R1456 vss.n131 vss.n130 0.0224072
R1457 vss.n142 vss.n138 0.0224072
R1458 vss.n144 vss.n142 0.0224072
R1459 vss.n148 vss.n144 0.0224072
R1460 vss.n150 vss.n148 0.0224072
R1461 vss.n154 vss.n150 0.0224072
R1462 vss.n156 vss.n154 0.0224072
R1463 vss.n160 vss.n156 0.0224072
R1464 vss.n162 vss.n160 0.0224072
R1465 vss.n166 vss.n162 0.0224072
R1466 vss.n168 vss.n166 0.0224072
R1467 vss.n172 vss.n168 0.0224072
R1468 vss.n174 vss.n172 0.0224072
R1469 vss.n671 vss.n667 0.0196441
R1470 vss.n762 vss.n757 0.0194732
R1471 vss.n415 vss.n412 0.0194732
R1472 vss.n349 vss.n345 0.0193053
R1473 vss.n695 vss.n694 0.018518
R1474 vss.n664 vss.n663 0.0176904
R1475 vss.n664 vss.n662 0.0176904
R1476 vss.n769 vss.n768 0.0176904
R1477 vss.n757 vss.n756 0.0176904
R1478 vss.n825 vss.n823 0.0176904
R1479 vss.n796 vss.n794 0.0176904
R1480 vss.n825 vss.n824 0.0176904
R1481 vss.n796 vss.n795 0.0176904
R1482 vss.n357 vss.n356 0.0176904
R1483 vss.n345 vss.n344 0.0176904
R1484 vss.n478 vss.n476 0.0176904
R1485 vss.n448 vss.n446 0.0176904
R1486 vss.n478 vss.n477 0.0176904
R1487 vss.n448 vss.n447 0.0176904
R1488 vss.n422 vss.n421 0.0176904
R1489 vss.n412 vss.n411 0.0176904
R1490 vss vss.n1002 0.0173269
R1491 vss.n754 vss.n749 0.016125
R1492 vss.n757 vss.n755 0.016125
R1493 vss.n409 vss.n404 0.016125
R1494 vss.n412 vss.n410 0.016125
R1495 vss.n342 vss.n337 0.0159867
R1496 vss.n345 vss.n343 0.0159867
R1497 vss.n694 vss.n692 0.0145766
R1498 vss.n49 vss.n43 0.0140309
R1499 vss.n137 vss.n131 0.0140309
R1500 vss.n665 vss.n664 0.0134505
R1501 vss.n770 vss.n769 0.0127768
R1502 vss.n423 vss.n422 0.0127768
R1503 vss.n358 vss.n357 0.0126681
R1504 vss.n691 vss.n686 0.0100721
R1505 vss.n686 vss.n682 0.0100721
R1506 vss.n682 vss.n680 0.0100721
R1507 vss.n680 vss.n678 0.0100721
R1508 vss.n678 vss.n674 0.0100721
R1509 vss.n733 vss.n729 0.0100721
R1510 vss.n735 vss.n733 0.0100721
R1511 vss.n705 vss.n700 0.0100721
R1512 vss.n720 vss.n717 0.0100721
R1513 vss.n321 vss.n319 0.0100721
R1514 vss.n319 vss.n314 0.0100721
R1515 vss.n388 vss.n384 0.0100721
R1516 vss.n390 vss.n388 0.0100721
R1517 vss.n767 vss.n762 0.00998661
R1518 vss.n769 vss.n767 0.00998661
R1519 vss.n777 vss.n774 0.00998661
R1520 vss.n790 vss.n786 0.00998661
R1521 vss.n420 vss.n415 0.00998661
R1522 vss.n422 vss.n420 0.00998661
R1523 vss.n430 vss.n427 0.00998661
R1524 vss.n442 vss.n439 0.00998661
R1525 vss.n355 vss.n349 0.00990266
R1526 vss.n357 vss.n355 0.00990266
R1527 vss.n365 vss.n362 0.00990266
R1528 vss.n380 vss.n376 0.00990266
R1529 vss.n721 vss.n720 0.00950901
R1530 vss.n791 vss.n790 0.00942857
R1531 vss.n443 vss.n442 0.00942857
R1532 vss.n381 vss.n380 0.00934956
R1533 vss.n50 vss.n49 0.00887629
R1534 vss.n138 vss.n137 0.00887629
R1535 vss.n652 vss.n651 0.00747072
R1536 vss.n651 vss.n650 0.00747072
R1537 vss.n700 vss.n696 0.00725676
R1538 vss.n774 vss.n770 0.00719643
R1539 vss.n427 vss.n423 0.00719643
R1540 vss.n362 vss.n358 0.00713717
R1541 vss.n833 vss.n825 0.00635399
R1542 vss.n486 vss.n478 0.00635399
R1543 vss.n667 vss.n665 0.00556757
R1544 vss.n692 vss.n691 0.00556757
R1545 vss.n792 vss.n721 0.00556757
R1546 vss.n792 vss.n791 0.00552232
R1547 vss.n444 vss.n443 0.00552232
R1548 vss.n444 vss.n381 0.00547788
R1549 vss.n834 vss.n833 0.00532094
R1550 vss.n487 vss.n486 0.00532094
R1551 vss.n825 vss.n822 0.00480441
R1552 vss.n478 vss.n475 0.00480441
R1553 vss.n871 vss.n835 0.00446006
R1554 vss.n521 vss.n488 0.00446006
R1555 vss.n696 vss.n695 0.00444144
R1556 vss.n755 vss.n735 0.00387838
R1557 vss.n410 vss.n390 0.00387838
R1558 vss.n755 vss.n754 0.00384821
R1559 vss.n410 vss.n409 0.00384821
R1560 vss.n343 vss.n342 0.00381858
R1561 vss.n811 vss.n796 0.003427
R1562 vss.n835 vss.n834 0.003427
R1563 vss.n464 vss.n448 0.003427
R1564 vss.n488 vss.n487 0.003427
R1565 vss.n724 vss.n722 0.00340353
R1566 vss.n311 vss.n309 0.00340353
R1567 vss.n821 vss.n813 0.00272259
R1568 vss.n474 vss.n466 0.00272259
R1569 vss.n710 vss.n708 0.00218919
R1570 vss.n782 vss.n780 0.00217411
R1571 vss.n435 vss.n433 0.00217411
R1572 vss.n370 vss.n368 0.00215929
R1573 vss.n871 vss.n843 0.00211903
R1574 vss.n521 vss.n500 0.00211903
R1575 vss.n822 vss.n821 0.00204959
R1576 vss.n475 vss.n474 0.00204959
R1577 vss.n813 vss.n811 0.00190551
R1578 vss.n466 vss.n464 0.00190551
R1579 vss.n793 vss.n792 0.00187741
R1580 vss.n445 vss.n444 0.00187741
R1581 vss.n664 vss.n652 0.00162613
R1582 vss.n695 vss.n671 0.00162613
R1583 vss.n343 vss.n321 0.00162613
R1584 vss.n872 vss.n871 0.00117218
R1585 vss.n522 vss.n521 0.00117218
R1586 vss.n210 vss.n209 0.00114971
R1587 vss.n276 vss.n275 0.00114971
R1588 vss.n969 vss.n968 0.00114971
R1589 vss.n909 vss.n908 0.00114971
R1590 vss.n619 vss.n618 0.00114971
R1591 vss.n558 vss.n557 0.00114971
R1592 vss.n726 vss.n724 0.00106306
R1593 vss.n311 vss.n308 0.00106306
R1594 vss.n49 vss.n48 0.00101178
R1595 vss.n137 vss.n136 0.00101178
R1596 vss.n813 vss.n812 0.00100251
R1597 vss.n466 vss.n465 0.00100251
R1598 vss.n872 vss.n649 0.00100144
R1599 vss.n522 vss.n306 0.00100144
R1600 vss.n796 vss.n793 0.000672176
R1601 vss.n448 vss.n445 0.000672176
R1602 vss.n708 vss.n706 0.000507886
R1603 vss.n780 vss.n778 0.000507886
R1604 vss.n433 vss.n431 0.000507886
R1605 vss.n368 vss.n366 0.000506749
R1606 vss.n710 vss.n709 0.000504067
R1607 vss.n782 vss.n781 0.000504067
R1608 vss.n435 vss.n434 0.000504067
R1609 vss.n370 vss.n369 0.000503481
R1610 vss.n724 vss.n723 0.000502566
R1611 vss.n311 vss.n310 0.000502566
R1612 vss.n726 vss.n725 0.000501438
R1613 vss.n308 vss.n307 0.000501438
R1614 vss.n708 vss.n707 0.000501244
R1615 vss.n780 vss.n779 0.000501244
R1616 vss.n368 vss.n367 0.000501244
R1617 vss.n433 vss.n432 0.000501244
R1618 a_n178_n2405.n2 a_n178_n2405.t14 68.4774
R1619 a_n178_n2405.n8 a_n178_n2405.t3 68.1157
R1620 a_n178_n2405.n6 a_n178_n2405.t7 67.9642
R1621 a_n178_n2405.n5 a_n178_n2405.t13 67.9642
R1622 a_n178_n2405.n4 a_n178_n2405.t15 67.9642
R1623 a_n178_n2405.n3 a_n178_n2405.t9 67.9642
R1624 a_n178_n2405.n2 a_n178_n2405.t12 67.9642
R1625 a_n178_n2405.n7 a_n178_n2405.t5 67.9642
R1626 a_n178_n2405.n18 a_n178_n2405.t1 17.4005
R1627 a_n178_n2405.n18 a_n178_n2405.t0 17.4005
R1628 a_n178_n2405.n10 a_n178_n2405.t2 17.4005
R1629 a_n178_n2405.n10 a_n178_n2405.t11 17.4005
R1630 a_n178_n2405.n13 a_n178_n2405.t8 5.7135
R1631 a_n178_n2405.n13 a_n178_n2405.t6 5.7135
R1632 a_n178_n2405.n21 a_n178_n2405.t4 5.7135
R1633 a_n178_n2405.t10 a_n178_n2405.n21 5.7135
R1634 a_n178_n2405.n14 a_n178_n2405.n13 1.21671
R1635 a_n178_n2405.n21 a_n178_n2405.n20 1.21671
R1636 a_n178_n2405.n9 a_n178_n2405.n2 0.633447
R1637 a_n178_n2405.n17 a_n178_n2405.n4 0.63175
R1638 a_n178_n2405.n1 a_n178_n2405.n11 0.555788
R1639 a_n178_n2405.n0 a_n178_n2405.n19 0.555788
R1640 a_n178_n2405.n4 a_n178_n2405.n16 0.550981
R1641 a_n178_n2405.n1 a_n178_n2405.n10 0.490863
R1642 a_n178_n2405.n0 a_n178_n2405.n18 0.488494
R1643 a_n178_n2405.n0 a_n178_n2405.n17 0.48175
R1644 a_n178_n2405.n1 a_n178_n2405.n9 0.48175
R1645 a_n178_n2405.n20 a_n178_n2405.n3 0.481269
R1646 a_n178_n2405.n6 a_n178_n2405.n14 0.481269
R1647 a_n178_n2405.n6 a_n178_n2405.n12 0.478282
R1648 a_n178_n2405.n4 a_n178_n2405.n15 0.478282
R1649 a_n178_n2405.n15 a_n178_n2405.n5 0.477583
R1650 a_n178_n2405.n12 a_n178_n2405.n7 0.477583
R1651 a_n178_n2405.n7 a_n178_n2405.n1 0.168596
R1652 a_n178_n2405.n3 a_n178_n2405.n0 0.168596
R1653 a_n178_n2405.n20 a_n178_n2405.n8 0.161036
R1654 a_n178_n2405.n5 a_n178_n2405.n6 1.26379
R1655 a_n3216_n2108.n17 a_n3216_n2108.n16 3175.18
R1656 a_n3216_n2108.n9 a_n3216_n2108.t3 18.9369
R1657 a_n3216_n2108.n9 a_n3216_n2108.t4 18.9346
R1658 a_n3216_n2108.n8 a_n3216_n2108.t2 18.8017
R1659 a_n3216_n2108.n8 a_n3216_n2108.t5 18.7979
R1660 a_n3216_n2108.n16 a_n3216_n2108.n0 9.3005
R1661 a_n3216_n2108.n16 a_n3216_n2108.n15 9.3005
R1662 a_n3216_n2108.n4 a_n3216_n2108.n1 9.10459
R1663 a_n3216_n2108.n11 a_n3216_n2108.n10 5.22377
R1664 a_n3216_n2108.n11 a_n3216_n2108.t0 4.99149
R1665 a_n3216_n2108.n4 a_n3216_n2108.n3 3.25237
R1666 a_n3216_n2108.n10 a_n3216_n2108.n8 2.57868
R1667 a_n3216_n2108.n12 a_n3216_n2108.n11 1.66518
R1668 a_n3216_n2108.n15 a_n3216_n2108.n14 1.30881
R1669 a_n3216_n2108.n10 a_n3216_n2108.n9 0.148227
R1670 a_n3216_n2108.n15 a_n3216_n2108.n4 0.0526884
R1671 a_n3216_n2108.n14 a_n3216_n2108.n13 0.0426677
R1672 a_n3216_n2108.n14 a_n3216_n2108.n7 0.0318735
R1673 a_n3216_n2108.n13 a_n3216_n2108.n12 0.016125
R1674 a_n3216_n2108.n7 a_n3216_n2108.n6 0.00577108
R1675 a_n3216_n2108.n6 a_n3216_n2108.n5 0.00263488
R1676 a_n3216_n2108.n3 a_n3216_n2108.n2 0.00117383
R1677 a_n3216_n2108.n2 a_n3216_n2108.t1 0.00101765
R1678 vtemp.n4 vtemp.t1 17.4005
R1679 vtemp.n4 vtemp.t2 17.4005
R1680 vtemp.n1 vtemp.t0 17.4005
R1681 vtemp.n1 vtemp.t3 17.4005
R1682 vtemp.n3 vtemp.t7 5.7135
R1683 vtemp.n3 vtemp.t5 5.7135
R1684 vtemp.n0 vtemp.t4 5.7135
R1685 vtemp.n0 vtemp.t6 5.7135
R1686 vtemp vtemp.n6 3.87576
R1687 vtemp.n6 vtemp.n5 2.56122
R1688 vtemp.n5 vtemp.n3 0.571731
R1689 vtemp.n2 vtemp.n0 0.569904
R1690 vtemp.n5 vtemp.n4 0.300087
R1691 vtemp.n2 vtemp.n1 0.300087
R1692 vtemp.n6 vtemp.n2 0.00352842
C0 a_n5752_n1958# a_n5810_n2748# 0.0726f
C1 vdd a_62_n3136# 0.0216f
C2 a_n5752_n2774# vdd 0.797f
C3 a_n5752_n1958# a_n5752_n3086# 1.38e-19
C4 a_n5752_n2774# a_n5810_n2748# 0.112f
C5 vdd vtemp 1.05f
C6 a_n5752_n2774# a_n5752_n3086# 0.324f
C7 a_n5752_n1958# a_n5752_n2774# 0.458f
C8 a_n5752_n2774# a_62_n3136# 1.46f
C9 a_n5810_n2748# vdd 0.132f
C10 vtemp a_62_n3136# 0.505f
C11 a_n5752_n3086# vdd 0.412f
C12 a_n5752_n2774# vtemp 0.00245f
C13 a_n5810_n2748# a_n5752_n3086# 0.0623f
C14 a_n5752_n1958# vdd 0.664f
.ends

