magic
tech sky130A
magscale 1 2
timestamp 1680390383
<< pwell >>
rect -307 -2008 307 2008
<< psubdiff >>
rect -271 1938 -175 1972
rect 175 1938 271 1972
rect -271 1876 -237 1938
rect 237 1876 271 1938
rect -271 -1938 -237 -1876
rect 237 -1938 271 -1876
rect -271 -1972 -175 -1938
rect 175 -1972 271 -1938
<< psubdiffcont >>
rect -175 1938 175 1972
rect -271 -1876 -237 1876
rect 237 -1876 271 1876
rect -175 -1972 175 -1938
<< xpolycontact >>
rect -141 1410 141 1842
rect -141 -1842 141 -1410
<< xpolyres >>
rect -141 -1410 141 1410
<< locali >>
rect -271 1938 -175 1972
rect 175 1938 271 1972
rect -271 1876 -237 1938
rect 237 1876 271 1938
rect -271 -1938 -237 -1876
rect 237 -1938 271 -1876
rect -271 -1972 -175 -1938
rect 175 -1972 271 -1938
<< viali >>
rect -125 1427 125 1824
rect -125 -1824 125 -1427
<< metal1 >>
rect -131 1824 131 1836
rect -131 1427 -125 1824
rect 125 1427 131 1824
rect -131 1415 131 1427
rect -131 -1427 131 -1415
rect -131 -1824 -125 -1427
rect 125 -1824 131 -1427
rect -131 -1836 131 -1824
<< res1p41 >>
rect -143 -1412 143 1412
<< properties >>
string FIXED_BBOX -254 -1955 254 1955
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 14.1 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 20.266k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
