* NGSPICE file created from ring_oscillator.ext - technology: sky130A

.subckt ring_oscillator vtemp vosc vss vdd
X0 a_2140_n4622.t0 vosc.t2 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=2e+06u
X1 vosc.t1 a_3744_n4622.t2 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=2e+06u
X2 a_2140_n4622.t1 vosc.t3 vss.t1 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3 vosc vtemp vss sky130_fd_pr__cap_var_lvt w=5e+06u l=5e+06u
X4 vosc.t0 a_3744_n4622.t3 vss.t5 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X5 a_3744_n4622.t0 a_2140_n4622.t3 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=2e+06u
X6 a_3744_n4622.t1 a_2140_n4622.t4 vss.t2 vss sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X7 a_2140_n4622.t0 vtemp vss sky130_fd_pr__cap_var_lvt w=5e+06u l=5e+06u
X8 a_3744_n4622.t0 vtemp vss sky130_fd_pr__cap_var_lvt w=5e+06u l=5e+06u
R0 vosc.n0 vosc.t2 152.33
R1 vosc.n0 vosc.t3 54.846
R2 vosc.n1 vosc.t4 14.094
R3 vosc.n3 vosc.n0 10.163
R4 vosc.n1 vosc.t0 4.35
R5 vosc.n2 vosc.t1 3.596
R6 vosc.n3 vosc.n2 0.732
R7 vosc.n2 vosc.n1 0.469
R8 vosc vosc.n3 0.342
R9 vdd.n17 vdd.t0 110.711
R10 vdd.n204 vdd.t2 110.711
R11 vdd.n391 vdd.t4 110.711
R12 vdd.n25 vdd.n22 12.923
R13 vdd.n212 vdd.n209 12.923
R14 vdd.n399 vdd.n396 12.923
R15 vdd.n185 vdd.n184 9.3
R16 vdd.n27 vdd.n26 9.3
R17 vdd.n30 vdd.n29 9.3
R18 vdd.n32 vdd.n31 9.3
R19 vdd.n35 vdd.n34 9.3
R20 vdd.n37 vdd.n36 9.3
R21 vdd.n40 vdd.n39 9.3
R22 vdd.n42 vdd.n41 9.3
R23 vdd.n45 vdd.n44 9.3
R24 vdd.n47 vdd.n46 9.3
R25 vdd.n50 vdd.n49 9.3
R26 vdd.n52 vdd.n51 9.3
R27 vdd.n55 vdd.n54 9.3
R28 vdd.n57 vdd.n56 9.3
R29 vdd.n60 vdd.n59 9.3
R30 vdd.n62 vdd.n61 9.3
R31 vdd.n65 vdd.n64 9.3
R32 vdd.n67 vdd.n66 9.3
R33 vdd.n70 vdd.n69 9.3
R34 vdd.n72 vdd.n71 9.3
R35 vdd.n75 vdd.n74 9.3
R36 vdd.n77 vdd.n76 9.3
R37 vdd.n80 vdd.n79 9.3
R38 vdd.n82 vdd.n81 9.3
R39 vdd.n85 vdd.n84 9.3
R40 vdd.n87 vdd.n86 9.3
R41 vdd.n90 vdd.n89 9.3
R42 vdd.n92 vdd.n91 9.3
R43 vdd.n95 vdd.n94 9.3
R44 vdd.n97 vdd.n96 9.3
R45 vdd.n100 vdd.n99 9.3
R46 vdd.n102 vdd.n101 9.3
R47 vdd.n105 vdd.n104 9.3
R48 vdd.n108 vdd.n107 9.3
R49 vdd.n110 vdd.n109 9.3
R50 vdd.n113 vdd.n112 9.3
R51 vdd.n115 vdd.n114 9.3
R52 vdd.n118 vdd.n117 9.3
R53 vdd.n120 vdd.n119 9.3
R54 vdd.n123 vdd.n122 9.3
R55 vdd.n125 vdd.n124 9.3
R56 vdd.n128 vdd.n127 9.3
R57 vdd.n130 vdd.n129 9.3
R58 vdd.n133 vdd.n132 9.3
R59 vdd.n135 vdd.n134 9.3
R60 vdd.n138 vdd.n137 9.3
R61 vdd.n140 vdd.n139 9.3
R62 vdd.n143 vdd.n142 9.3
R63 vdd.n145 vdd.n144 9.3
R64 vdd.n148 vdd.n147 9.3
R65 vdd.n150 vdd.n149 9.3
R66 vdd.n153 vdd.n152 9.3
R67 vdd.n155 vdd.n154 9.3
R68 vdd.n158 vdd.n157 9.3
R69 vdd.n160 vdd.n159 9.3
R70 vdd.n163 vdd.n162 9.3
R71 vdd.n165 vdd.n164 9.3
R72 vdd.n168 vdd.n167 9.3
R73 vdd.n170 vdd.n169 9.3
R74 vdd.n173 vdd.n172 9.3
R75 vdd.n175 vdd.n174 9.3
R76 vdd.n178 vdd.n177 9.3
R77 vdd.n180 vdd.n179 9.3
R78 vdd.n183 vdd.n182 9.3
R79 vdd.n214 vdd.n213 9.3
R80 vdd.n217 vdd.n216 9.3
R81 vdd.n219 vdd.n218 9.3
R82 vdd.n222 vdd.n221 9.3
R83 vdd.n224 vdd.n223 9.3
R84 vdd.n227 vdd.n226 9.3
R85 vdd.n229 vdd.n228 9.3
R86 vdd.n232 vdd.n231 9.3
R87 vdd.n234 vdd.n233 9.3
R88 vdd.n237 vdd.n236 9.3
R89 vdd.n239 vdd.n238 9.3
R90 vdd.n242 vdd.n241 9.3
R91 vdd.n244 vdd.n243 9.3
R92 vdd.n247 vdd.n246 9.3
R93 vdd.n249 vdd.n248 9.3
R94 vdd.n252 vdd.n251 9.3
R95 vdd.n254 vdd.n253 9.3
R96 vdd.n257 vdd.n256 9.3
R97 vdd.n259 vdd.n258 9.3
R98 vdd.n262 vdd.n261 9.3
R99 vdd.n264 vdd.n263 9.3
R100 vdd.n267 vdd.n266 9.3
R101 vdd.n269 vdd.n268 9.3
R102 vdd.n272 vdd.n271 9.3
R103 vdd.n274 vdd.n273 9.3
R104 vdd.n277 vdd.n276 9.3
R105 vdd.n279 vdd.n278 9.3
R106 vdd.n282 vdd.n281 9.3
R107 vdd.n284 vdd.n283 9.3
R108 vdd.n287 vdd.n286 9.3
R109 vdd.n289 vdd.n288 9.3
R110 vdd.n292 vdd.n291 9.3
R111 vdd.n295 vdd.n294 9.3
R112 vdd.n297 vdd.n296 9.3
R113 vdd.n300 vdd.n299 9.3
R114 vdd.n302 vdd.n301 9.3
R115 vdd.n305 vdd.n304 9.3
R116 vdd.n307 vdd.n306 9.3
R117 vdd.n310 vdd.n309 9.3
R118 vdd.n312 vdd.n311 9.3
R119 vdd.n315 vdd.n314 9.3
R120 vdd.n317 vdd.n316 9.3
R121 vdd.n320 vdd.n319 9.3
R122 vdd.n322 vdd.n321 9.3
R123 vdd.n325 vdd.n324 9.3
R124 vdd.n327 vdd.n326 9.3
R125 vdd.n330 vdd.n329 9.3
R126 vdd.n332 vdd.n331 9.3
R127 vdd.n335 vdd.n334 9.3
R128 vdd.n337 vdd.n336 9.3
R129 vdd.n340 vdd.n339 9.3
R130 vdd.n342 vdd.n341 9.3
R131 vdd.n345 vdd.n344 9.3
R132 vdd.n347 vdd.n346 9.3
R133 vdd.n350 vdd.n349 9.3
R134 vdd.n352 vdd.n351 9.3
R135 vdd.n355 vdd.n354 9.3
R136 vdd.n357 vdd.n356 9.3
R137 vdd.n360 vdd.n359 9.3
R138 vdd.n362 vdd.n361 9.3
R139 vdd.n365 vdd.n364 9.3
R140 vdd.n367 vdd.n366 9.3
R141 vdd.n370 vdd.n369 9.3
R142 vdd.n372 vdd.n371 9.3
R143 vdd.n401 vdd.n400 9.3
R144 vdd.n404 vdd.n403 9.3
R145 vdd.n406 vdd.n405 9.3
R146 vdd.n409 vdd.n408 9.3
R147 vdd.n411 vdd.n410 9.3
R148 vdd.n414 vdd.n413 9.3
R149 vdd.n416 vdd.n415 9.3
R150 vdd.n419 vdd.n418 9.3
R151 vdd.n421 vdd.n420 9.3
R152 vdd.n424 vdd.n423 9.3
R153 vdd.n426 vdd.n425 9.3
R154 vdd.n429 vdd.n428 9.3
R155 vdd.n431 vdd.n430 9.3
R156 vdd.n434 vdd.n433 9.3
R157 vdd.n436 vdd.n435 9.3
R158 vdd.n439 vdd.n438 9.3
R159 vdd.n441 vdd.n440 9.3
R160 vdd.n444 vdd.n443 9.3
R161 vdd.n446 vdd.n445 9.3
R162 vdd.n449 vdd.n448 9.3
R163 vdd.n451 vdd.n450 9.3
R164 vdd.n454 vdd.n453 9.3
R165 vdd.n456 vdd.n455 9.3
R166 vdd.n459 vdd.n458 9.3
R167 vdd.n461 vdd.n460 9.3
R168 vdd.n464 vdd.n463 9.3
R169 vdd.n466 vdd.n465 9.3
R170 vdd.n469 vdd.n468 9.3
R171 vdd.n471 vdd.n470 9.3
R172 vdd.n474 vdd.n473 9.3
R173 vdd.n476 vdd.n475 9.3
R174 vdd.n479 vdd.n478 9.3
R175 vdd.n482 vdd.n481 9.3
R176 vdd.n484 vdd.n483 9.3
R177 vdd.n487 vdd.n486 9.3
R178 vdd.n489 vdd.n488 9.3
R179 vdd.n492 vdd.n491 9.3
R180 vdd.n494 vdd.n493 9.3
R181 vdd.n497 vdd.n496 9.3
R182 vdd.n499 vdd.n498 9.3
R183 vdd.n502 vdd.n501 9.3
R184 vdd.n504 vdd.n503 9.3
R185 vdd.n507 vdd.n506 9.3
R186 vdd.n509 vdd.n508 9.3
R187 vdd.n512 vdd.n511 9.3
R188 vdd.n514 vdd.n513 9.3
R189 vdd.n517 vdd.n516 9.3
R190 vdd.n519 vdd.n518 9.3
R191 vdd.n522 vdd.n521 9.3
R192 vdd.n524 vdd.n523 9.3
R193 vdd.n527 vdd.n526 9.3
R194 vdd.n529 vdd.n528 9.3
R195 vdd.n532 vdd.n531 9.3
R196 vdd.n534 vdd.n533 9.3
R197 vdd.n537 vdd.n536 9.3
R198 vdd.n539 vdd.n538 9.3
R199 vdd.n542 vdd.n541 9.3
R200 vdd.n544 vdd.n543 9.3
R201 vdd.n547 vdd.n546 9.3
R202 vdd.n549 vdd.n548 9.3
R203 vdd.n552 vdd.n551 9.3
R204 vdd.n554 vdd.n553 9.3
R205 vdd.n557 vdd.n556 9.3
R206 vdd.n559 vdd.n558 9.3
R207 vdd.n24 vdd.n23 8.855
R208 vdd.n29 vdd.n28 8.855
R209 vdd.n34 vdd.n33 8.855
R210 vdd.n39 vdd.n38 8.855
R211 vdd.n44 vdd.n43 8.855
R212 vdd.n49 vdd.n48 8.855
R213 vdd.n54 vdd.n53 8.855
R214 vdd.n59 vdd.n58 8.855
R215 vdd.n64 vdd.n63 8.855
R216 vdd.n69 vdd.n68 8.855
R217 vdd.n74 vdd.n73 8.855
R218 vdd.n79 vdd.n78 8.855
R219 vdd.n84 vdd.n83 8.855
R220 vdd.n89 vdd.n88 8.855
R221 vdd.n94 vdd.n93 8.855
R222 vdd.n99 vdd.n98 8.855
R223 vdd.n20 vdd.n19 8.855
R224 vdd.n107 vdd.n106 8.855
R225 vdd.n112 vdd.n111 8.855
R226 vdd.n117 vdd.n116 8.855
R227 vdd.n122 vdd.n121 8.855
R228 vdd.n127 vdd.n126 8.855
R229 vdd.n132 vdd.n131 8.855
R230 vdd.n137 vdd.n136 8.855
R231 vdd.n142 vdd.n141 8.855
R232 vdd.n147 vdd.n146 8.855
R233 vdd.n152 vdd.n151 8.855
R234 vdd.n157 vdd.n156 8.855
R235 vdd.n162 vdd.n161 8.855
R236 vdd.n167 vdd.n166 8.855
R237 vdd.n172 vdd.n171 8.855
R238 vdd.n177 vdd.n176 8.855
R239 vdd.n182 vdd.n181 8.855
R240 vdd.n211 vdd.n210 8.855
R241 vdd.n216 vdd.n215 8.855
R242 vdd.n221 vdd.n220 8.855
R243 vdd.n226 vdd.n225 8.855
R244 vdd.n231 vdd.n230 8.855
R245 vdd.n236 vdd.n235 8.855
R246 vdd.n241 vdd.n240 8.855
R247 vdd.n246 vdd.n245 8.855
R248 vdd.n251 vdd.n250 8.855
R249 vdd.n256 vdd.n255 8.855
R250 vdd.n261 vdd.n260 8.855
R251 vdd.n266 vdd.n265 8.855
R252 vdd.n271 vdd.n270 8.855
R253 vdd.n276 vdd.n275 8.855
R254 vdd.n281 vdd.n280 8.855
R255 vdd.n286 vdd.n285 8.855
R256 vdd.n207 vdd.n206 8.855
R257 vdd.n294 vdd.n293 8.855
R258 vdd.n299 vdd.n298 8.855
R259 vdd.n304 vdd.n303 8.855
R260 vdd.n309 vdd.n308 8.855
R261 vdd.n314 vdd.n313 8.855
R262 vdd.n319 vdd.n318 8.855
R263 vdd.n324 vdd.n323 8.855
R264 vdd.n329 vdd.n328 8.855
R265 vdd.n334 vdd.n333 8.855
R266 vdd.n339 vdd.n338 8.855
R267 vdd.n344 vdd.n343 8.855
R268 vdd.n349 vdd.n348 8.855
R269 vdd.n354 vdd.n353 8.855
R270 vdd.n359 vdd.n358 8.855
R271 vdd.n364 vdd.n363 8.855
R272 vdd.n369 vdd.n368 8.855
R273 vdd.n398 vdd.n397 8.855
R274 vdd.n403 vdd.n402 8.855
R275 vdd.n408 vdd.n407 8.855
R276 vdd.n413 vdd.n412 8.855
R277 vdd.n418 vdd.n417 8.855
R278 vdd.n423 vdd.n422 8.855
R279 vdd.n428 vdd.n427 8.855
R280 vdd.n433 vdd.n432 8.855
R281 vdd.n438 vdd.n437 8.855
R282 vdd.n443 vdd.n442 8.855
R283 vdd.n448 vdd.n447 8.855
R284 vdd.n453 vdd.n452 8.855
R285 vdd.n458 vdd.n457 8.855
R286 vdd.n463 vdd.n462 8.855
R287 vdd.n468 vdd.n467 8.855
R288 vdd.n473 vdd.n472 8.855
R289 vdd.n394 vdd.n393 8.855
R290 vdd.n481 vdd.n480 8.855
R291 vdd.n486 vdd.n485 8.855
R292 vdd.n491 vdd.n490 8.855
R293 vdd.n496 vdd.n495 8.855
R294 vdd.n501 vdd.n500 8.855
R295 vdd.n506 vdd.n505 8.855
R296 vdd.n511 vdd.n510 8.855
R297 vdd.n516 vdd.n515 8.855
R298 vdd.n521 vdd.n520 8.855
R299 vdd.n526 vdd.n525 8.855
R300 vdd.n531 vdd.n530 8.855
R301 vdd.n536 vdd.n535 8.855
R302 vdd.n541 vdd.n540 8.855
R303 vdd.n546 vdd.n545 8.855
R304 vdd.n551 vdd.n550 8.855
R305 vdd.n556 vdd.n555 8.855
R306 vdd.n19 vdd.n18 7.775
R307 vdd.n206 vdd.n205 7.775
R308 vdd.n393 vdd.n392 7.775
R309 vdd.n186 vdd.n0 6.166
R310 vdd.n373 vdd.n187 6.166
R311 vdd.n560 vdd.n374 6.166
R312 vdd.n25 vdd.n24 5.571
R313 vdd.n212 vdd.n211 5.571
R314 vdd.n399 vdd.n398 5.571
R315 vdd.n103 vdd.t1 2.38
R316 vdd.n290 vdd.t3 2.38
R317 vdd.n477 vdd.t5 2.38
R318 vdd.n561 vdd.n560 0.783
R319 vdd.n27 vdd.n25 0.713
R320 vdd.n214 vdd.n212 0.713
R321 vdd.n401 vdd.n399 0.713
R322 vdd.n17 vdd.n16 0.54
R323 vdd.n17 vdd.n15 0.54
R324 vdd.n17 vdd.n14 0.54
R325 vdd.n17 vdd.n13 0.54
R326 vdd.n17 vdd.n12 0.54
R327 vdd.n17 vdd.n11 0.54
R328 vdd.n17 vdd.n10 0.54
R329 vdd.n17 vdd.n9 0.54
R330 vdd.n18 vdd.n17 0.54
R331 vdd.n17 vdd.n8 0.54
R332 vdd.n17 vdd.n7 0.54
R333 vdd.n17 vdd.n6 0.54
R334 vdd.n17 vdd.n5 0.54
R335 vdd.n17 vdd.n4 0.54
R336 vdd.n17 vdd.n3 0.54
R337 vdd.n17 vdd.n2 0.54
R338 vdd.n17 vdd.n1 0.54
R339 vdd.n204 vdd.n203 0.54
R340 vdd.n204 vdd.n202 0.54
R341 vdd.n204 vdd.n201 0.54
R342 vdd.n204 vdd.n200 0.54
R343 vdd.n204 vdd.n199 0.54
R344 vdd.n204 vdd.n198 0.54
R345 vdd.n204 vdd.n197 0.54
R346 vdd.n204 vdd.n196 0.54
R347 vdd.n205 vdd.n204 0.54
R348 vdd.n204 vdd.n195 0.54
R349 vdd.n204 vdd.n194 0.54
R350 vdd.n204 vdd.n193 0.54
R351 vdd.n204 vdd.n192 0.54
R352 vdd.n204 vdd.n191 0.54
R353 vdd.n204 vdd.n190 0.54
R354 vdd.n204 vdd.n189 0.54
R355 vdd.n204 vdd.n188 0.54
R356 vdd.n391 vdd.n390 0.54
R357 vdd.n391 vdd.n389 0.54
R358 vdd.n391 vdd.n388 0.54
R359 vdd.n391 vdd.n387 0.54
R360 vdd.n391 vdd.n386 0.54
R361 vdd.n391 vdd.n385 0.54
R362 vdd.n391 vdd.n384 0.54
R363 vdd.n391 vdd.n383 0.54
R364 vdd.n392 vdd.n391 0.54
R365 vdd.n391 vdd.n382 0.54
R366 vdd.n391 vdd.n381 0.54
R367 vdd.n391 vdd.n380 0.54
R368 vdd.n391 vdd.n379 0.54
R369 vdd.n391 vdd.n378 0.54
R370 vdd.n391 vdd.n377 0.54
R371 vdd.n391 vdd.n376 0.54
R372 vdd.n391 vdd.n375 0.54
R373 vdd.n562 vdd.n561 0.433
R374 vdd.n21 vdd.n20 0.362
R375 vdd.n208 vdd.n207 0.362
R376 vdd.n395 vdd.n394 0.362
R377 vdd.n562 vdd.n186 0.35
R378 vdd.n561 vdd.n373 0.35
R379 vdd vdd.n562 0.123
R380 vdd.n186 vdd.n185 0.039
R381 vdd.n373 vdd.n372 0.039
R382 vdd.n560 vdd.n559 0.039
R383 vdd.n185 vdd.n183 0.031
R384 vdd.n183 vdd.n180 0.031
R385 vdd.n180 vdd.n178 0.031
R386 vdd.n178 vdd.n175 0.031
R387 vdd.n175 vdd.n173 0.031
R388 vdd.n173 vdd.n170 0.031
R389 vdd.n170 vdd.n168 0.031
R390 vdd.n168 vdd.n165 0.031
R391 vdd.n165 vdd.n163 0.031
R392 vdd.n163 vdd.n160 0.031
R393 vdd.n160 vdd.n158 0.031
R394 vdd.n158 vdd.n155 0.031
R395 vdd.n155 vdd.n153 0.031
R396 vdd.n153 vdd.n150 0.031
R397 vdd.n150 vdd.n148 0.031
R398 vdd.n148 vdd.n145 0.031
R399 vdd.n145 vdd.n143 0.031
R400 vdd.n143 vdd.n140 0.031
R401 vdd.n140 vdd.n138 0.031
R402 vdd.n138 vdd.n135 0.031
R403 vdd.n135 vdd.n133 0.031
R404 vdd.n133 vdd.n130 0.031
R405 vdd.n130 vdd.n128 0.031
R406 vdd.n128 vdd.n125 0.031
R407 vdd.n125 vdd.n123 0.031
R408 vdd.n123 vdd.n120 0.031
R409 vdd.n120 vdd.n118 0.031
R410 vdd.n118 vdd.n115 0.031
R411 vdd.n115 vdd.n113 0.031
R412 vdd.n113 vdd.n110 0.031
R413 vdd.n110 vdd.n108 0.031
R414 vdd.n108 vdd.n105 0.031
R415 vdd.n105 vdd.n103 0.031
R416 vdd.n102 vdd.n100 0.031
R417 vdd.n100 vdd.n97 0.031
R418 vdd.n97 vdd.n95 0.031
R419 vdd.n95 vdd.n92 0.031
R420 vdd.n92 vdd.n90 0.031
R421 vdd.n90 vdd.n87 0.031
R422 vdd.n87 vdd.n85 0.031
R423 vdd.n85 vdd.n82 0.031
R424 vdd.n82 vdd.n80 0.031
R425 vdd.n80 vdd.n77 0.031
R426 vdd.n77 vdd.n75 0.031
R427 vdd.n75 vdd.n72 0.031
R428 vdd.n72 vdd.n70 0.031
R429 vdd.n70 vdd.n67 0.031
R430 vdd.n67 vdd.n65 0.031
R431 vdd.n65 vdd.n62 0.031
R432 vdd.n62 vdd.n60 0.031
R433 vdd.n60 vdd.n57 0.031
R434 vdd.n57 vdd.n55 0.031
R435 vdd.n55 vdd.n52 0.031
R436 vdd.n52 vdd.n50 0.031
R437 vdd.n50 vdd.n47 0.031
R438 vdd.n47 vdd.n45 0.031
R439 vdd.n45 vdd.n42 0.031
R440 vdd.n42 vdd.n40 0.031
R441 vdd.n40 vdd.n37 0.031
R442 vdd.n37 vdd.n35 0.031
R443 vdd.n35 vdd.n32 0.031
R444 vdd.n32 vdd.n30 0.031
R445 vdd.n30 vdd.n27 0.031
R446 vdd.n372 vdd.n370 0.031
R447 vdd.n370 vdd.n367 0.031
R448 vdd.n367 vdd.n365 0.031
R449 vdd.n365 vdd.n362 0.031
R450 vdd.n362 vdd.n360 0.031
R451 vdd.n360 vdd.n357 0.031
R452 vdd.n357 vdd.n355 0.031
R453 vdd.n355 vdd.n352 0.031
R454 vdd.n352 vdd.n350 0.031
R455 vdd.n350 vdd.n347 0.031
R456 vdd.n347 vdd.n345 0.031
R457 vdd.n345 vdd.n342 0.031
R458 vdd.n342 vdd.n340 0.031
R459 vdd.n340 vdd.n337 0.031
R460 vdd.n337 vdd.n335 0.031
R461 vdd.n335 vdd.n332 0.031
R462 vdd.n332 vdd.n330 0.031
R463 vdd.n330 vdd.n327 0.031
R464 vdd.n327 vdd.n325 0.031
R465 vdd.n325 vdd.n322 0.031
R466 vdd.n322 vdd.n320 0.031
R467 vdd.n320 vdd.n317 0.031
R468 vdd.n317 vdd.n315 0.031
R469 vdd.n315 vdd.n312 0.031
R470 vdd.n312 vdd.n310 0.031
R471 vdd.n310 vdd.n307 0.031
R472 vdd.n307 vdd.n305 0.031
R473 vdd.n305 vdd.n302 0.031
R474 vdd.n302 vdd.n300 0.031
R475 vdd.n300 vdd.n297 0.031
R476 vdd.n297 vdd.n295 0.031
R477 vdd.n295 vdd.n292 0.031
R478 vdd.n292 vdd.n290 0.031
R479 vdd.n289 vdd.n287 0.031
R480 vdd.n287 vdd.n284 0.031
R481 vdd.n284 vdd.n282 0.031
R482 vdd.n282 vdd.n279 0.031
R483 vdd.n279 vdd.n277 0.031
R484 vdd.n277 vdd.n274 0.031
R485 vdd.n274 vdd.n272 0.031
R486 vdd.n272 vdd.n269 0.031
R487 vdd.n269 vdd.n267 0.031
R488 vdd.n267 vdd.n264 0.031
R489 vdd.n264 vdd.n262 0.031
R490 vdd.n262 vdd.n259 0.031
R491 vdd.n259 vdd.n257 0.031
R492 vdd.n257 vdd.n254 0.031
R493 vdd.n254 vdd.n252 0.031
R494 vdd.n252 vdd.n249 0.031
R495 vdd.n249 vdd.n247 0.031
R496 vdd.n247 vdd.n244 0.031
R497 vdd.n244 vdd.n242 0.031
R498 vdd.n242 vdd.n239 0.031
R499 vdd.n239 vdd.n237 0.031
R500 vdd.n237 vdd.n234 0.031
R501 vdd.n234 vdd.n232 0.031
R502 vdd.n232 vdd.n229 0.031
R503 vdd.n229 vdd.n227 0.031
R504 vdd.n227 vdd.n224 0.031
R505 vdd.n224 vdd.n222 0.031
R506 vdd.n222 vdd.n219 0.031
R507 vdd.n219 vdd.n217 0.031
R508 vdd.n217 vdd.n214 0.031
R509 vdd.n559 vdd.n557 0.031
R510 vdd.n557 vdd.n554 0.031
R511 vdd.n554 vdd.n552 0.031
R512 vdd.n552 vdd.n549 0.031
R513 vdd.n549 vdd.n547 0.031
R514 vdd.n547 vdd.n544 0.031
R515 vdd.n544 vdd.n542 0.031
R516 vdd.n542 vdd.n539 0.031
R517 vdd.n539 vdd.n537 0.031
R518 vdd.n537 vdd.n534 0.031
R519 vdd.n534 vdd.n532 0.031
R520 vdd.n532 vdd.n529 0.031
R521 vdd.n529 vdd.n527 0.031
R522 vdd.n527 vdd.n524 0.031
R523 vdd.n524 vdd.n522 0.031
R524 vdd.n522 vdd.n519 0.031
R525 vdd.n519 vdd.n517 0.031
R526 vdd.n517 vdd.n514 0.031
R527 vdd.n514 vdd.n512 0.031
R528 vdd.n512 vdd.n509 0.031
R529 vdd.n509 vdd.n507 0.031
R530 vdd.n507 vdd.n504 0.031
R531 vdd.n504 vdd.n502 0.031
R532 vdd.n502 vdd.n499 0.031
R533 vdd.n499 vdd.n497 0.031
R534 vdd.n497 vdd.n494 0.031
R535 vdd.n494 vdd.n492 0.031
R536 vdd.n492 vdd.n489 0.031
R537 vdd.n489 vdd.n487 0.031
R538 vdd.n487 vdd.n484 0.031
R539 vdd.n484 vdd.n482 0.031
R540 vdd.n482 vdd.n479 0.031
R541 vdd.n479 vdd.n477 0.031
R542 vdd.n476 vdd.n474 0.031
R543 vdd.n474 vdd.n471 0.031
R544 vdd.n471 vdd.n469 0.031
R545 vdd.n469 vdd.n466 0.031
R546 vdd.n466 vdd.n464 0.031
R547 vdd.n464 vdd.n461 0.031
R548 vdd.n461 vdd.n459 0.031
R549 vdd.n459 vdd.n456 0.031
R550 vdd.n456 vdd.n454 0.031
R551 vdd.n454 vdd.n451 0.031
R552 vdd.n451 vdd.n449 0.031
R553 vdd.n449 vdd.n446 0.031
R554 vdd.n446 vdd.n444 0.031
R555 vdd.n444 vdd.n441 0.031
R556 vdd.n441 vdd.n439 0.031
R557 vdd.n439 vdd.n436 0.031
R558 vdd.n436 vdd.n434 0.031
R559 vdd.n434 vdd.n431 0.031
R560 vdd.n431 vdd.n429 0.031
R561 vdd.n429 vdd.n426 0.031
R562 vdd.n426 vdd.n424 0.031
R563 vdd.n424 vdd.n421 0.031
R564 vdd.n421 vdd.n419 0.031
R565 vdd.n419 vdd.n416 0.031
R566 vdd.n416 vdd.n414 0.031
R567 vdd.n414 vdd.n411 0.031
R568 vdd.n411 vdd.n409 0.031
R569 vdd.n409 vdd.n406 0.031
R570 vdd.n406 vdd.n404 0.031
R571 vdd.n404 vdd.n401 0.031
R572 vdd.n103 vdd.n102 0.03
R573 vdd.n290 vdd.n289 0.03
R574 vdd.n477 vdd.n476 0.03
R575 vdd.n103 vdd.n21 0.001
R576 vdd.n290 vdd.n208 0.001
R577 vdd.n477 vdd.n395 0.001
R578 a_2140_n4622.n0 a_2140_n4622.t3 152.33
R579 a_2140_n4622.n0 a_2140_n4622.t4 54.846
R580 a_2140_n4622.n1 a_2140_n4622.t2 14.096
R581 a_2140_n4622.n1 a_2140_n4622.n0 9.319
R582 a_2140_n4622.n2 a_2140_n4622.t1 4.35
R583 a_2140_n4622.t0 a_2140_n4622.n2 4.117
R584 a_2140_n4622.n2 a_2140_n4622.n1 0.22
R585 a_3744_n4622.n0 a_3744_n4622.t2 152.313
R586 a_3744_n4622.n0 a_3744_n4622.t3 54.829
R587 a_3744_n4622.n1 a_3744_n4622.t4 13.865
R588 a_3744_n4622.n1 a_3744_n4622.n0 9.317
R589 a_3744_n4622.n2 a_3744_n4622.t1 4.35
R590 a_3744_n4622.t0 a_3744_n4622.n2 4.117
R591 a_3744_n4622.n2 a_3744_n4622.n1 0.22
R592 vss.n211 vss.n210 9.3
R593 vss.n209 vss.n208 9.3
R594 vss.n206 vss.n205 9.3
R595 vss.n204 vss.n203 9.3
R596 vss.n201 vss.n200 9.3
R597 vss.n199 vss.n198 9.3
R598 vss.n196 vss.n195 9.3
R599 vss.n194 vss.n193 9.3
R600 vss.n191 vss.n190 9.3
R601 vss.n273 vss.n272 9.3
R602 vss.n271 vss.n270 9.3
R603 vss.n268 vss.n267 9.3
R604 vss.n266 vss.n265 9.3
R605 vss.n263 vss.n262 9.3
R606 vss.n261 vss.n260 9.3
R607 vss.n258 vss.n257 9.3
R608 vss.n256 vss.n255 9.3
R609 vss.n253 vss.n252 9.3
R610 vss.n251 vss.n250 9.3
R611 vss.n248 vss.n247 9.3
R612 vss.n242 vss.n241 9.3
R613 vss.n240 vss.n239 9.3
R614 vss.n237 vss.n236 9.3
R615 vss.n235 vss.n234 9.3
R616 vss.n232 vss.n231 9.3
R617 vss.n230 vss.n229 9.3
R618 vss.n227 vss.n226 9.3
R619 vss.n225 vss.n224 9.3
R620 vss.n222 vss.n221 9.3
R621 vss.n220 vss.n219 9.3
R622 vss.n217 vss.n216 9.3
R623 vss.n275 vss.n274 9.3
R624 vss.n119 vss.n118 9.3
R625 vss.n117 vss.n116 9.3
R626 vss.n114 vss.n113 9.3
R627 vss.n112 vss.n111 9.3
R628 vss.n109 vss.n108 9.3
R629 vss.n107 vss.n106 9.3
R630 vss.n104 vss.n103 9.3
R631 vss.n102 vss.n101 9.3
R632 vss.n99 vss.n98 9.3
R633 vss.n181 vss.n180 9.3
R634 vss.n179 vss.n178 9.3
R635 vss.n176 vss.n175 9.3
R636 vss.n174 vss.n173 9.3
R637 vss.n171 vss.n170 9.3
R638 vss.n169 vss.n168 9.3
R639 vss.n166 vss.n165 9.3
R640 vss.n164 vss.n163 9.3
R641 vss.n161 vss.n160 9.3
R642 vss.n159 vss.n158 9.3
R643 vss.n156 vss.n155 9.3
R644 vss.n150 vss.n149 9.3
R645 vss.n148 vss.n147 9.3
R646 vss.n145 vss.n144 9.3
R647 vss.n143 vss.n142 9.3
R648 vss.n140 vss.n139 9.3
R649 vss.n138 vss.n137 9.3
R650 vss.n135 vss.n134 9.3
R651 vss.n133 vss.n132 9.3
R652 vss.n130 vss.n129 9.3
R653 vss.n128 vss.n127 9.3
R654 vss.n125 vss.n124 9.3
R655 vss.n183 vss.n182 9.3
R656 vss.n27 vss.n26 9.3
R657 vss.n25 vss.n24 9.3
R658 vss.n22 vss.n21 9.3
R659 vss.n20 vss.n19 9.3
R660 vss.n17 vss.n16 9.3
R661 vss.n15 vss.n14 9.3
R662 vss.n12 vss.n11 9.3
R663 vss.n10 vss.n9 9.3
R664 vss.n7 vss.n6 9.3
R665 vss.n89 vss.n88 9.3
R666 vss.n87 vss.n86 9.3
R667 vss.n84 vss.n83 9.3
R668 vss.n82 vss.n81 9.3
R669 vss.n79 vss.n78 9.3
R670 vss.n77 vss.n76 9.3
R671 vss.n74 vss.n73 9.3
R672 vss.n72 vss.n71 9.3
R673 vss.n69 vss.n68 9.3
R674 vss.n67 vss.n66 9.3
R675 vss.n64 vss.n63 9.3
R676 vss.n58 vss.n57 9.3
R677 vss.n56 vss.n55 9.3
R678 vss.n53 vss.n52 9.3
R679 vss.n51 vss.n50 9.3
R680 vss.n48 vss.n47 9.3
R681 vss.n46 vss.n45 9.3
R682 vss.n43 vss.n42 9.3
R683 vss.n41 vss.n40 9.3
R684 vss.n38 vss.n37 9.3
R685 vss.n36 vss.n35 9.3
R686 vss.n33 vss.n32 9.3
R687 vss.n91 vss.n90 9.3
R688 vss.n270 vss.n269 9.154
R689 vss.n208 vss.n207 9.154
R690 vss.n203 vss.n202 9.154
R691 vss.n198 vss.n197 9.154
R692 vss.n193 vss.n192 9.154
R693 vss.n187 vss.n186 9.154
R694 vss.n265 vss.n264 9.154
R695 vss.n260 vss.n259 9.154
R696 vss.n255 vss.n254 9.154
R697 vss.n250 vss.n249 9.154
R698 vss.n185 vss.n184 9.154
R699 vss.n244 vss.n243 9.154
R700 vss.n239 vss.n238 9.154
R701 vss.n234 vss.n233 9.154
R702 vss.n229 vss.n228 9.154
R703 vss.n224 vss.n223 9.154
R704 vss.n219 vss.n218 9.154
R705 vss.n178 vss.n177 9.154
R706 vss.n116 vss.n115 9.154
R707 vss.n111 vss.n110 9.154
R708 vss.n106 vss.n105 9.154
R709 vss.n101 vss.n100 9.154
R710 vss.n95 vss.n94 9.154
R711 vss.n173 vss.n172 9.154
R712 vss.n168 vss.n167 9.154
R713 vss.n163 vss.n162 9.154
R714 vss.n158 vss.n157 9.154
R715 vss.n93 vss.n92 9.154
R716 vss.n152 vss.n151 9.154
R717 vss.n147 vss.n146 9.154
R718 vss.n142 vss.n141 9.154
R719 vss.n137 vss.n136 9.154
R720 vss.n132 vss.n131 9.154
R721 vss.n127 vss.n126 9.154
R722 vss.n86 vss.n85 9.154
R723 vss.n24 vss.n23 9.154
R724 vss.n19 vss.n18 9.154
R725 vss.n14 vss.n13 9.154
R726 vss.n9 vss.n8 9.154
R727 vss.n3 vss.n2 9.154
R728 vss.n81 vss.n80 9.154
R729 vss.n76 vss.n75 9.154
R730 vss.n71 vss.n70 9.154
R731 vss.n66 vss.n65 9.154
R732 vss.n1 vss.n0 9.154
R733 vss.n60 vss.n59 9.154
R734 vss.n55 vss.n54 9.154
R735 vss.n50 vss.n49 9.154
R736 vss.n45 vss.n44 9.154
R737 vss.n40 vss.n39 9.154
R738 vss.n35 vss.n34 9.154
R739 vss.n215 vss.n214 6.539
R740 vss.n123 vss.n122 6.539
R741 vss.n31 vss.n30 6.539
R742 vss.n213 vss.n212 6.209
R743 vss.n121 vss.n120 6.209
R744 vss.n29 vss.n28 6.209
R745 vss.n246 vss.n185 5.949
R746 vss.n154 vss.n93 5.949
R747 vss.n62 vss.n1 5.949
R748 vss.n188 vss.t1 4.35
R749 vss.n96 vss.t2 4.35
R750 vss.n4 vss.t5 4.35
R751 vss.n245 vss.n244 3.787
R752 vss.n153 vss.n152 3.787
R753 vss.n61 vss.n60 3.787
R754 vss.n189 vss.n187 3.512
R755 vss.n97 vss.n95 3.512
R756 vss.n5 vss.n3 3.512
R757 vss vss.n91 0.67
R758 vss.n277 vss.n276 0.434
R759 vss.n277 vss.n183 0.404
R760 vss.n276 vss.n275 0.402
R761 vss.n123 vss.n121 0.329
R762 vss.n215 vss.n213 0.327
R763 vss.n31 vss.n29 0.327
R764 vss vss.n277 0.164
R765 vss.n276 vss 0.107
R766 vss.n248 vss.n246 0.053
R767 vss.n156 vss.n154 0.053
R768 vss.n64 vss.n62 0.053
R769 vss.n217 vss.n215 0.047
R770 vss.n245 vss.n242 0.047
R771 vss.n125 vss.n123 0.047
R772 vss.n153 vss.n150 0.047
R773 vss.n33 vss.n31 0.047
R774 vss.n61 vss.n58 0.047
R775 vss.n246 vss.n245 0.046
R776 vss.n154 vss.n153 0.046
R777 vss.n62 vss.n61 0.046
R778 vss.n220 vss.n217 0.036
R779 vss.n222 vss.n220 0.036
R780 vss.n225 vss.n222 0.036
R781 vss.n227 vss.n225 0.036
R782 vss.n230 vss.n227 0.036
R783 vss.n232 vss.n230 0.036
R784 vss.n235 vss.n232 0.036
R785 vss.n237 vss.n235 0.036
R786 vss.n240 vss.n237 0.036
R787 vss.n242 vss.n240 0.036
R788 vss.n251 vss.n248 0.036
R789 vss.n253 vss.n251 0.036
R790 vss.n256 vss.n253 0.036
R791 vss.n258 vss.n256 0.036
R792 vss.n261 vss.n258 0.036
R793 vss.n263 vss.n261 0.036
R794 vss.n266 vss.n263 0.036
R795 vss.n268 vss.n266 0.036
R796 vss.n271 vss.n268 0.036
R797 vss.n273 vss.n271 0.036
R798 vss.n275 vss.n273 0.036
R799 vss.n128 vss.n125 0.036
R800 vss.n130 vss.n128 0.036
R801 vss.n133 vss.n130 0.036
R802 vss.n135 vss.n133 0.036
R803 vss.n138 vss.n135 0.036
R804 vss.n140 vss.n138 0.036
R805 vss.n143 vss.n140 0.036
R806 vss.n145 vss.n143 0.036
R807 vss.n148 vss.n145 0.036
R808 vss.n150 vss.n148 0.036
R809 vss.n159 vss.n156 0.036
R810 vss.n161 vss.n159 0.036
R811 vss.n164 vss.n161 0.036
R812 vss.n166 vss.n164 0.036
R813 vss.n169 vss.n166 0.036
R814 vss.n171 vss.n169 0.036
R815 vss.n174 vss.n171 0.036
R816 vss.n176 vss.n174 0.036
R817 vss.n179 vss.n176 0.036
R818 vss.n181 vss.n179 0.036
R819 vss.n183 vss.n181 0.036
R820 vss.n36 vss.n33 0.036
R821 vss.n38 vss.n36 0.036
R822 vss.n41 vss.n38 0.036
R823 vss.n43 vss.n41 0.036
R824 vss.n46 vss.n43 0.036
R825 vss.n48 vss.n46 0.036
R826 vss.n51 vss.n48 0.036
R827 vss.n53 vss.n51 0.036
R828 vss.n56 vss.n53 0.036
R829 vss.n58 vss.n56 0.036
R830 vss.n67 vss.n64 0.036
R831 vss.n69 vss.n67 0.036
R832 vss.n72 vss.n69 0.036
R833 vss.n74 vss.n72 0.036
R834 vss.n77 vss.n74 0.036
R835 vss.n79 vss.n77 0.036
R836 vss.n82 vss.n79 0.036
R837 vss.n84 vss.n82 0.036
R838 vss.n87 vss.n84 0.036
R839 vss.n89 vss.n87 0.036
R840 vss.n91 vss.n89 0.036
R841 vss.n191 vss.n189 0.028
R842 vss.n99 vss.n97 0.028
R843 vss.n7 vss.n5 0.028
R844 vss.n213 vss.n211 0.028
R845 vss.n121 vss.n119 0.028
R846 vss.n29 vss.n27 0.028
R847 vss.n194 vss.n191 0.022
R848 vss.n196 vss.n194 0.022
R849 vss.n199 vss.n196 0.022
R850 vss.n201 vss.n199 0.022
R851 vss.n204 vss.n201 0.022
R852 vss.n206 vss.n204 0.022
R853 vss.n209 vss.n206 0.022
R854 vss.n211 vss.n209 0.022
R855 vss.n102 vss.n99 0.022
R856 vss.n104 vss.n102 0.022
R857 vss.n107 vss.n104 0.022
R858 vss.n109 vss.n107 0.022
R859 vss.n112 vss.n109 0.022
R860 vss.n114 vss.n112 0.022
R861 vss.n117 vss.n114 0.022
R862 vss.n119 vss.n117 0.022
R863 vss.n10 vss.n7 0.022
R864 vss.n12 vss.n10 0.022
R865 vss.n15 vss.n12 0.022
R866 vss.n17 vss.n15 0.022
R867 vss.n20 vss.n17 0.022
R868 vss.n22 vss.n20 0.022
R869 vss.n25 vss.n22 0.022
R870 vss.n27 vss.n25 0.022
R871 vss.n189 vss.n188 0.004
R872 vss.n97 vss.n96 0.004
R873 vss.n5 vss.n4 0.004
R874 vtemp.n1 vtemp.t1 8.087
R875 vtemp.n0 vtemp.t2 8.087
R876 vtemp.n0 vtemp.t0 9.059
R877 vtemp vtemp.n1 1.082
R878 vtemp.n1 vtemp.n0 0.963
C0 vdd vosc 1.65fF
C1 vdd vtemp 0.07fF
C2 vtemp vosc 6.73fF
.ends

