magic
tech sky130A
magscale 1 2
timestamp 1680262531
<< nwell >>
rect -396 -619 396 619
<< pmoslvt >>
rect -200 -400 200 400
<< pdiff >>
rect -258 388 -200 400
rect -258 -388 -246 388
rect -212 -388 -200 388
rect -258 -400 -200 -388
rect 200 388 258 400
rect 200 -388 212 388
rect 246 -388 258 388
rect 200 -400 258 -388
<< pdiffc >>
rect -246 -388 -212 388
rect 212 -388 246 388
<< nsubdiff >>
rect -360 549 -264 583
rect 264 549 360 583
rect -360 487 -326 549
rect 326 487 360 549
rect -360 -549 -326 -487
rect 326 -549 360 -487
rect -360 -583 -264 -549
rect 264 -583 360 -549
<< nsubdiffcont >>
rect -264 549 264 583
rect -360 -487 -326 487
rect 326 -487 360 487
rect -264 -583 264 -549
<< poly >>
rect -200 481 200 497
rect -200 447 -184 481
rect 184 447 200 481
rect -200 400 200 447
rect -200 -447 200 -400
rect -200 -481 -184 -447
rect 184 -481 200 -447
rect -200 -497 200 -481
<< polycont >>
rect -184 447 184 481
rect -184 -481 184 -447
<< locali >>
rect -360 549 -264 583
rect 264 549 360 583
rect -360 487 -326 549
rect 326 487 360 549
rect -200 447 -184 481
rect 184 447 200 481
rect -246 388 -212 404
rect -246 -404 -212 -388
rect 212 388 246 404
rect 212 -404 246 -388
rect -200 -481 -184 -447
rect 184 -481 200 -447
rect -360 -549 -326 -487
rect 326 -549 360 -487
rect -360 -583 -264 -549
rect 264 -583 360 -549
<< viali >>
rect -184 447 184 481
rect -246 -388 -212 388
rect 212 -388 246 388
rect -184 -481 184 -447
<< metal1 >>
rect -196 481 196 487
rect -196 447 -184 481
rect 184 447 196 481
rect -196 441 196 447
rect -252 388 -206 400
rect -252 -388 -246 388
rect -212 -388 -206 388
rect -252 -400 -206 -388
rect 206 388 252 400
rect 206 -388 212 388
rect 246 -388 252 388
rect 206 -400 252 -388
rect -196 -447 196 -441
rect -196 -481 -184 -447
rect 184 -481 196 -447
rect -196 -487 196 -481
<< properties >>
string FIXED_BBOX -343 -566 343 566
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
