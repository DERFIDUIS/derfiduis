magic
tech sky130A
magscale 1 2
timestamp 1681063793
<< nwell >>
rect 12354 -3060 12420 -1860
rect 12758 -3060 12872 -1860
rect 13162 -3060 13276 -1860
rect 13566 -3060 13680 -1860
rect 13970 -3060 14084 -1860
rect 14374 -3060 14488 -1860
rect 14826 -3060 14892 -1860
<< ndiff >>
rect 12658 -4436 12660 -3436
rect 12906 -4436 12908 -3436
rect 12994 -4436 12996 -3436
rect 13242 -4436 13244 -3436
rect 13330 -4436 13332 -3436
rect 13578 -4436 13580 -3436
rect 13666 -4436 13668 -3436
rect 13914 -4436 13916 -3436
rect 14002 -4436 14004 -3436
rect 14250 -4436 14252 -3436
rect 14338 -4436 14340 -3436
rect 14586 -4436 14588 -3436
<< pdiff >>
rect 12454 -2960 12456 -1960
rect 12770 -2960 12772 -1960
rect 12858 -2960 12860 -1960
rect 13174 -2960 13176 -1960
rect 13262 -2960 13264 -1960
rect 13578 -2960 13580 -1960
rect 13666 -2960 13668 -1960
rect 13982 -2960 13984 -1960
rect 14070 -2960 14072 -1960
rect 14386 -2960 14388 -1960
rect 14474 -2960 14476 -1960
rect 14790 -2960 14792 -1960
<< psubdiff >>
rect 12594 -3490 12658 -3436
rect 12594 -3524 12598 -3490
rect 12632 -3524 12658 -3490
rect 12594 -3558 12658 -3524
rect 12594 -3592 12598 -3558
rect 12632 -3592 12658 -3558
rect 12594 -3626 12658 -3592
rect 12594 -3660 12598 -3626
rect 12632 -3660 12658 -3626
rect 12594 -3694 12658 -3660
rect 12594 -3728 12598 -3694
rect 12632 -3728 12658 -3694
rect 12594 -3762 12658 -3728
rect 12594 -3796 12598 -3762
rect 12632 -3796 12658 -3762
rect 12594 -3830 12658 -3796
rect 12594 -3864 12598 -3830
rect 12632 -3864 12658 -3830
rect 12594 -3898 12658 -3864
rect 12594 -3932 12598 -3898
rect 12632 -3932 12658 -3898
rect 12594 -3966 12658 -3932
rect 12594 -4000 12598 -3966
rect 12632 -4000 12658 -3966
rect 12594 -4034 12658 -4000
rect 12594 -4068 12598 -4034
rect 12632 -4068 12658 -4034
rect 12594 -4102 12658 -4068
rect 12594 -4136 12598 -4102
rect 12632 -4136 12658 -4102
rect 12594 -4170 12658 -4136
rect 12594 -4204 12598 -4170
rect 12632 -4204 12658 -4170
rect 12594 -4238 12658 -4204
rect 12594 -4272 12598 -4238
rect 12632 -4272 12658 -4238
rect 12594 -4306 12658 -4272
rect 12594 -4340 12598 -4306
rect 12632 -4340 12658 -4306
rect 12594 -4374 12658 -4340
rect 12594 -4408 12598 -4374
rect 12632 -4408 12658 -4374
rect 12594 -4436 12658 -4408
rect 12908 -3464 12994 -3436
rect 12908 -3498 12934 -3464
rect 12968 -3498 12994 -3464
rect 12908 -3532 12994 -3498
rect 12908 -3566 12934 -3532
rect 12968 -3566 12994 -3532
rect 12908 -3600 12994 -3566
rect 12908 -3634 12934 -3600
rect 12968 -3634 12994 -3600
rect 12908 -3668 12994 -3634
rect 12908 -3702 12934 -3668
rect 12968 -3702 12994 -3668
rect 12908 -3736 12994 -3702
rect 12908 -3770 12934 -3736
rect 12968 -3770 12994 -3736
rect 12908 -3804 12994 -3770
rect 12908 -3838 12934 -3804
rect 12968 -3838 12994 -3804
rect 12908 -3872 12994 -3838
rect 12908 -3906 12934 -3872
rect 12968 -3906 12994 -3872
rect 12908 -3940 12994 -3906
rect 12908 -3974 12934 -3940
rect 12968 -3974 12994 -3940
rect 12908 -4008 12994 -3974
rect 12908 -4042 12934 -4008
rect 12968 -4042 12994 -4008
rect 12908 -4076 12994 -4042
rect 12908 -4110 12934 -4076
rect 12968 -4110 12994 -4076
rect 12908 -4144 12994 -4110
rect 12908 -4178 12934 -4144
rect 12968 -4178 12994 -4144
rect 12908 -4212 12994 -4178
rect 12908 -4246 12934 -4212
rect 12968 -4246 12994 -4212
rect 12908 -4280 12994 -4246
rect 12908 -4314 12934 -4280
rect 12968 -4314 12994 -4280
rect 12908 -4348 12994 -4314
rect 12908 -4382 12934 -4348
rect 12968 -4382 12994 -4348
rect 12908 -4436 12994 -4382
rect 13244 -3464 13330 -3436
rect 13244 -3498 13270 -3464
rect 13304 -3498 13330 -3464
rect 13244 -3532 13330 -3498
rect 13244 -3566 13270 -3532
rect 13304 -3566 13330 -3532
rect 13244 -3600 13330 -3566
rect 13244 -3634 13270 -3600
rect 13304 -3634 13330 -3600
rect 13244 -3668 13330 -3634
rect 13244 -3702 13270 -3668
rect 13304 -3702 13330 -3668
rect 13244 -3736 13330 -3702
rect 13244 -3770 13270 -3736
rect 13304 -3770 13330 -3736
rect 13244 -3804 13330 -3770
rect 13244 -3838 13270 -3804
rect 13304 -3838 13330 -3804
rect 13244 -3872 13330 -3838
rect 13244 -3906 13270 -3872
rect 13304 -3906 13330 -3872
rect 13244 -3940 13330 -3906
rect 13244 -3974 13270 -3940
rect 13304 -3974 13330 -3940
rect 13244 -4008 13330 -3974
rect 13244 -4042 13270 -4008
rect 13304 -4042 13330 -4008
rect 13244 -4076 13330 -4042
rect 13244 -4110 13270 -4076
rect 13304 -4110 13330 -4076
rect 13244 -4144 13330 -4110
rect 13244 -4178 13270 -4144
rect 13304 -4178 13330 -4144
rect 13244 -4212 13330 -4178
rect 13244 -4246 13270 -4212
rect 13304 -4246 13330 -4212
rect 13244 -4280 13330 -4246
rect 13244 -4314 13270 -4280
rect 13304 -4314 13330 -4280
rect 13244 -4348 13330 -4314
rect 13244 -4382 13270 -4348
rect 13304 -4382 13330 -4348
rect 13244 -4436 13330 -4382
rect 13580 -3464 13666 -3436
rect 13580 -3498 13606 -3464
rect 13640 -3498 13666 -3464
rect 13580 -3532 13666 -3498
rect 13580 -3566 13606 -3532
rect 13640 -3566 13666 -3532
rect 13580 -3600 13666 -3566
rect 13580 -3634 13606 -3600
rect 13640 -3634 13666 -3600
rect 13580 -3668 13666 -3634
rect 13580 -3702 13606 -3668
rect 13640 -3702 13666 -3668
rect 13580 -3736 13666 -3702
rect 13580 -3770 13606 -3736
rect 13640 -3770 13666 -3736
rect 13580 -3804 13666 -3770
rect 13580 -3838 13606 -3804
rect 13640 -3838 13666 -3804
rect 13580 -3872 13666 -3838
rect 13580 -3906 13606 -3872
rect 13640 -3906 13666 -3872
rect 13580 -3940 13666 -3906
rect 13580 -3974 13606 -3940
rect 13640 -3974 13666 -3940
rect 13580 -4008 13666 -3974
rect 13580 -4042 13606 -4008
rect 13640 -4042 13666 -4008
rect 13580 -4076 13666 -4042
rect 13580 -4110 13606 -4076
rect 13640 -4110 13666 -4076
rect 13580 -4144 13666 -4110
rect 13580 -4178 13606 -4144
rect 13640 -4178 13666 -4144
rect 13580 -4212 13666 -4178
rect 13580 -4246 13606 -4212
rect 13640 -4246 13666 -4212
rect 13580 -4280 13666 -4246
rect 13580 -4314 13606 -4280
rect 13640 -4314 13666 -4280
rect 13580 -4348 13666 -4314
rect 13580 -4382 13606 -4348
rect 13640 -4382 13666 -4348
rect 13580 -4436 13666 -4382
rect 13916 -3464 14002 -3436
rect 13916 -3498 13942 -3464
rect 13976 -3498 14002 -3464
rect 13916 -3532 14002 -3498
rect 13916 -3566 13942 -3532
rect 13976 -3566 14002 -3532
rect 13916 -3600 14002 -3566
rect 13916 -3634 13942 -3600
rect 13976 -3634 14002 -3600
rect 13916 -3668 14002 -3634
rect 13916 -3702 13942 -3668
rect 13976 -3702 14002 -3668
rect 13916 -3736 14002 -3702
rect 13916 -3770 13942 -3736
rect 13976 -3770 14002 -3736
rect 13916 -3804 14002 -3770
rect 13916 -3838 13942 -3804
rect 13976 -3838 14002 -3804
rect 13916 -3872 14002 -3838
rect 13916 -3906 13942 -3872
rect 13976 -3906 14002 -3872
rect 13916 -3940 14002 -3906
rect 13916 -3974 13942 -3940
rect 13976 -3974 14002 -3940
rect 13916 -4008 14002 -3974
rect 13916 -4042 13942 -4008
rect 13976 -4042 14002 -4008
rect 13916 -4076 14002 -4042
rect 13916 -4110 13942 -4076
rect 13976 -4110 14002 -4076
rect 13916 -4144 14002 -4110
rect 13916 -4178 13942 -4144
rect 13976 -4178 14002 -4144
rect 13916 -4212 14002 -4178
rect 13916 -4246 13942 -4212
rect 13976 -4246 14002 -4212
rect 13916 -4280 14002 -4246
rect 13916 -4314 13942 -4280
rect 13976 -4314 14002 -4280
rect 13916 -4348 14002 -4314
rect 13916 -4382 13942 -4348
rect 13976 -4382 14002 -4348
rect 13916 -4436 14002 -4382
rect 14252 -3464 14338 -3436
rect 14252 -3498 14278 -3464
rect 14312 -3498 14338 -3464
rect 14252 -3532 14338 -3498
rect 14252 -3566 14278 -3532
rect 14312 -3566 14338 -3532
rect 14252 -3600 14338 -3566
rect 14252 -3634 14278 -3600
rect 14312 -3634 14338 -3600
rect 14252 -3668 14338 -3634
rect 14252 -3702 14278 -3668
rect 14312 -3702 14338 -3668
rect 14252 -3736 14338 -3702
rect 14252 -3770 14278 -3736
rect 14312 -3770 14338 -3736
rect 14252 -3804 14338 -3770
rect 14252 -3838 14278 -3804
rect 14312 -3838 14338 -3804
rect 14252 -3872 14338 -3838
rect 14252 -3906 14278 -3872
rect 14312 -3906 14338 -3872
rect 14252 -3940 14338 -3906
rect 14252 -3974 14278 -3940
rect 14312 -3974 14338 -3940
rect 14252 -4008 14338 -3974
rect 14252 -4042 14278 -4008
rect 14312 -4042 14338 -4008
rect 14252 -4076 14338 -4042
rect 14252 -4110 14278 -4076
rect 14312 -4110 14338 -4076
rect 14252 -4144 14338 -4110
rect 14252 -4178 14278 -4144
rect 14312 -4178 14338 -4144
rect 14252 -4212 14338 -4178
rect 14252 -4246 14278 -4212
rect 14312 -4246 14338 -4212
rect 14252 -4280 14338 -4246
rect 14252 -4314 14278 -4280
rect 14312 -4314 14338 -4280
rect 14252 -4348 14338 -4314
rect 14252 -4382 14278 -4348
rect 14312 -4382 14338 -4348
rect 14252 -4436 14338 -4382
rect 14588 -3464 14652 -3436
rect 14588 -3498 14614 -3464
rect 14648 -3498 14652 -3464
rect 14588 -3532 14652 -3498
rect 14588 -3566 14614 -3532
rect 14648 -3566 14652 -3532
rect 14588 -3600 14652 -3566
rect 14588 -3634 14614 -3600
rect 14648 -3634 14652 -3600
rect 14588 -3668 14652 -3634
rect 14588 -3702 14614 -3668
rect 14648 -3702 14652 -3668
rect 14588 -3736 14652 -3702
rect 14588 -3770 14614 -3736
rect 14648 -3770 14652 -3736
rect 14588 -3804 14652 -3770
rect 14588 -3838 14614 -3804
rect 14648 -3838 14652 -3804
rect 14588 -3872 14652 -3838
rect 14588 -3906 14614 -3872
rect 14648 -3906 14652 -3872
rect 14588 -3940 14652 -3906
rect 14588 -3974 14614 -3940
rect 14648 -3974 14652 -3940
rect 14588 -4008 14652 -3974
rect 14588 -4042 14614 -4008
rect 14648 -4042 14652 -4008
rect 14588 -4076 14652 -4042
rect 14588 -4110 14614 -4076
rect 14648 -4110 14652 -4076
rect 14588 -4144 14652 -4110
rect 14588 -4178 14614 -4144
rect 14648 -4178 14652 -4144
rect 14588 -4212 14652 -4178
rect 14588 -4246 14614 -4212
rect 14648 -4246 14652 -4212
rect 14588 -4280 14652 -4246
rect 14588 -4314 14614 -4280
rect 14648 -4314 14652 -4280
rect 14588 -4348 14652 -4314
rect 14588 -4382 14614 -4348
rect 14648 -4382 14652 -4348
rect 14588 -4436 14652 -4382
<< nsubdiff >>
rect 12390 -2014 12454 -1960
rect 12390 -2048 12394 -2014
rect 12428 -2048 12454 -2014
rect 12390 -2082 12454 -2048
rect 12390 -2116 12394 -2082
rect 12428 -2116 12454 -2082
rect 12390 -2150 12454 -2116
rect 12390 -2184 12394 -2150
rect 12428 -2184 12454 -2150
rect 12390 -2218 12454 -2184
rect 12390 -2252 12394 -2218
rect 12428 -2252 12454 -2218
rect 12390 -2286 12454 -2252
rect 12390 -2320 12394 -2286
rect 12428 -2320 12454 -2286
rect 12390 -2354 12454 -2320
rect 12390 -2388 12394 -2354
rect 12428 -2388 12454 -2354
rect 12390 -2422 12454 -2388
rect 12390 -2456 12394 -2422
rect 12428 -2456 12454 -2422
rect 12390 -2490 12454 -2456
rect 12390 -2524 12394 -2490
rect 12428 -2524 12454 -2490
rect 12390 -2558 12454 -2524
rect 12390 -2592 12394 -2558
rect 12428 -2592 12454 -2558
rect 12390 -2626 12454 -2592
rect 12390 -2660 12394 -2626
rect 12428 -2660 12454 -2626
rect 12390 -2694 12454 -2660
rect 12390 -2728 12394 -2694
rect 12428 -2728 12454 -2694
rect 12390 -2762 12454 -2728
rect 12390 -2796 12394 -2762
rect 12428 -2796 12454 -2762
rect 12390 -2830 12454 -2796
rect 12390 -2864 12394 -2830
rect 12428 -2864 12454 -2830
rect 12390 -2898 12454 -2864
rect 12390 -2932 12394 -2898
rect 12428 -2932 12454 -2898
rect 12390 -2960 12454 -2932
rect 12772 -1988 12858 -1960
rect 12772 -2022 12798 -1988
rect 12832 -2022 12858 -1988
rect 12772 -2056 12858 -2022
rect 12772 -2090 12798 -2056
rect 12832 -2090 12858 -2056
rect 12772 -2124 12858 -2090
rect 12772 -2158 12798 -2124
rect 12832 -2158 12858 -2124
rect 12772 -2192 12858 -2158
rect 12772 -2226 12798 -2192
rect 12832 -2226 12858 -2192
rect 12772 -2260 12858 -2226
rect 12772 -2294 12798 -2260
rect 12832 -2294 12858 -2260
rect 12772 -2328 12858 -2294
rect 12772 -2362 12798 -2328
rect 12832 -2362 12858 -2328
rect 12772 -2396 12858 -2362
rect 12772 -2430 12798 -2396
rect 12832 -2430 12858 -2396
rect 12772 -2464 12858 -2430
rect 12772 -2498 12798 -2464
rect 12832 -2498 12858 -2464
rect 12772 -2532 12858 -2498
rect 12772 -2566 12798 -2532
rect 12832 -2566 12858 -2532
rect 12772 -2600 12858 -2566
rect 12772 -2634 12798 -2600
rect 12832 -2634 12858 -2600
rect 12772 -2668 12858 -2634
rect 12772 -2702 12798 -2668
rect 12832 -2702 12858 -2668
rect 12772 -2736 12858 -2702
rect 12772 -2770 12798 -2736
rect 12832 -2770 12858 -2736
rect 12772 -2804 12858 -2770
rect 12772 -2838 12798 -2804
rect 12832 -2838 12858 -2804
rect 12772 -2872 12858 -2838
rect 12772 -2906 12798 -2872
rect 12832 -2906 12858 -2872
rect 12772 -2960 12858 -2906
rect 13176 -1988 13262 -1960
rect 13176 -2022 13202 -1988
rect 13236 -2022 13262 -1988
rect 13176 -2056 13262 -2022
rect 13176 -2090 13202 -2056
rect 13236 -2090 13262 -2056
rect 13176 -2124 13262 -2090
rect 13176 -2158 13202 -2124
rect 13236 -2158 13262 -2124
rect 13176 -2192 13262 -2158
rect 13176 -2226 13202 -2192
rect 13236 -2226 13262 -2192
rect 13176 -2260 13262 -2226
rect 13176 -2294 13202 -2260
rect 13236 -2294 13262 -2260
rect 13176 -2328 13262 -2294
rect 13176 -2362 13202 -2328
rect 13236 -2362 13262 -2328
rect 13176 -2396 13262 -2362
rect 13176 -2430 13202 -2396
rect 13236 -2430 13262 -2396
rect 13176 -2464 13262 -2430
rect 13176 -2498 13202 -2464
rect 13236 -2498 13262 -2464
rect 13176 -2532 13262 -2498
rect 13176 -2566 13202 -2532
rect 13236 -2566 13262 -2532
rect 13176 -2600 13262 -2566
rect 13176 -2634 13202 -2600
rect 13236 -2634 13262 -2600
rect 13176 -2668 13262 -2634
rect 13176 -2702 13202 -2668
rect 13236 -2702 13262 -2668
rect 13176 -2736 13262 -2702
rect 13176 -2770 13202 -2736
rect 13236 -2770 13262 -2736
rect 13176 -2804 13262 -2770
rect 13176 -2838 13202 -2804
rect 13236 -2838 13262 -2804
rect 13176 -2872 13262 -2838
rect 13176 -2906 13202 -2872
rect 13236 -2906 13262 -2872
rect 13176 -2960 13262 -2906
rect 13580 -1988 13666 -1960
rect 13580 -2022 13606 -1988
rect 13640 -2022 13666 -1988
rect 13580 -2056 13666 -2022
rect 13580 -2090 13606 -2056
rect 13640 -2090 13666 -2056
rect 13580 -2124 13666 -2090
rect 13580 -2158 13606 -2124
rect 13640 -2158 13666 -2124
rect 13580 -2192 13666 -2158
rect 13580 -2226 13606 -2192
rect 13640 -2226 13666 -2192
rect 13580 -2260 13666 -2226
rect 13580 -2294 13606 -2260
rect 13640 -2294 13666 -2260
rect 13580 -2328 13666 -2294
rect 13580 -2362 13606 -2328
rect 13640 -2362 13666 -2328
rect 13580 -2396 13666 -2362
rect 13580 -2430 13606 -2396
rect 13640 -2430 13666 -2396
rect 13580 -2464 13666 -2430
rect 13580 -2498 13606 -2464
rect 13640 -2498 13666 -2464
rect 13580 -2532 13666 -2498
rect 13580 -2566 13606 -2532
rect 13640 -2566 13666 -2532
rect 13580 -2600 13666 -2566
rect 13580 -2634 13606 -2600
rect 13640 -2634 13666 -2600
rect 13580 -2668 13666 -2634
rect 13580 -2702 13606 -2668
rect 13640 -2702 13666 -2668
rect 13580 -2736 13666 -2702
rect 13580 -2770 13606 -2736
rect 13640 -2770 13666 -2736
rect 13580 -2804 13666 -2770
rect 13580 -2838 13606 -2804
rect 13640 -2838 13666 -2804
rect 13580 -2872 13666 -2838
rect 13580 -2906 13606 -2872
rect 13640 -2906 13666 -2872
rect 13580 -2960 13666 -2906
rect 13984 -1988 14070 -1960
rect 13984 -2022 14010 -1988
rect 14044 -2022 14070 -1988
rect 13984 -2056 14070 -2022
rect 13984 -2090 14010 -2056
rect 14044 -2090 14070 -2056
rect 13984 -2124 14070 -2090
rect 13984 -2158 14010 -2124
rect 14044 -2158 14070 -2124
rect 13984 -2192 14070 -2158
rect 13984 -2226 14010 -2192
rect 14044 -2226 14070 -2192
rect 13984 -2260 14070 -2226
rect 13984 -2294 14010 -2260
rect 14044 -2294 14070 -2260
rect 13984 -2328 14070 -2294
rect 13984 -2362 14010 -2328
rect 14044 -2362 14070 -2328
rect 13984 -2396 14070 -2362
rect 13984 -2430 14010 -2396
rect 14044 -2430 14070 -2396
rect 13984 -2464 14070 -2430
rect 13984 -2498 14010 -2464
rect 14044 -2498 14070 -2464
rect 13984 -2532 14070 -2498
rect 13984 -2566 14010 -2532
rect 14044 -2566 14070 -2532
rect 13984 -2600 14070 -2566
rect 13984 -2634 14010 -2600
rect 14044 -2634 14070 -2600
rect 13984 -2668 14070 -2634
rect 13984 -2702 14010 -2668
rect 14044 -2702 14070 -2668
rect 13984 -2736 14070 -2702
rect 13984 -2770 14010 -2736
rect 14044 -2770 14070 -2736
rect 13984 -2804 14070 -2770
rect 13984 -2838 14010 -2804
rect 14044 -2838 14070 -2804
rect 13984 -2872 14070 -2838
rect 13984 -2906 14010 -2872
rect 14044 -2906 14070 -2872
rect 13984 -2960 14070 -2906
rect 14388 -1988 14474 -1960
rect 14388 -2022 14414 -1988
rect 14448 -2022 14474 -1988
rect 14388 -2056 14474 -2022
rect 14388 -2090 14414 -2056
rect 14448 -2090 14474 -2056
rect 14388 -2124 14474 -2090
rect 14388 -2158 14414 -2124
rect 14448 -2158 14474 -2124
rect 14388 -2192 14474 -2158
rect 14388 -2226 14414 -2192
rect 14448 -2226 14474 -2192
rect 14388 -2260 14474 -2226
rect 14388 -2294 14414 -2260
rect 14448 -2294 14474 -2260
rect 14388 -2328 14474 -2294
rect 14388 -2362 14414 -2328
rect 14448 -2362 14474 -2328
rect 14388 -2396 14474 -2362
rect 14388 -2430 14414 -2396
rect 14448 -2430 14474 -2396
rect 14388 -2464 14474 -2430
rect 14388 -2498 14414 -2464
rect 14448 -2498 14474 -2464
rect 14388 -2532 14474 -2498
rect 14388 -2566 14414 -2532
rect 14448 -2566 14474 -2532
rect 14388 -2600 14474 -2566
rect 14388 -2634 14414 -2600
rect 14448 -2634 14474 -2600
rect 14388 -2668 14474 -2634
rect 14388 -2702 14414 -2668
rect 14448 -2702 14474 -2668
rect 14388 -2736 14474 -2702
rect 14388 -2770 14414 -2736
rect 14448 -2770 14474 -2736
rect 14388 -2804 14474 -2770
rect 14388 -2838 14414 -2804
rect 14448 -2838 14474 -2804
rect 14388 -2872 14474 -2838
rect 14388 -2906 14414 -2872
rect 14448 -2906 14474 -2872
rect 14388 -2960 14474 -2906
rect 14792 -1988 14856 -1960
rect 14792 -2022 14818 -1988
rect 14852 -2022 14856 -1988
rect 14792 -2056 14856 -2022
rect 14792 -2090 14818 -2056
rect 14852 -2090 14856 -2056
rect 14792 -2124 14856 -2090
rect 14792 -2158 14818 -2124
rect 14852 -2158 14856 -2124
rect 14792 -2192 14856 -2158
rect 14792 -2226 14818 -2192
rect 14852 -2226 14856 -2192
rect 14792 -2260 14856 -2226
rect 14792 -2294 14818 -2260
rect 14852 -2294 14856 -2260
rect 14792 -2328 14856 -2294
rect 14792 -2362 14818 -2328
rect 14852 -2362 14856 -2328
rect 14792 -2396 14856 -2362
rect 14792 -2430 14818 -2396
rect 14852 -2430 14856 -2396
rect 14792 -2464 14856 -2430
rect 14792 -2498 14818 -2464
rect 14852 -2498 14856 -2464
rect 14792 -2532 14856 -2498
rect 14792 -2566 14818 -2532
rect 14852 -2566 14856 -2532
rect 14792 -2600 14856 -2566
rect 14792 -2634 14818 -2600
rect 14852 -2634 14856 -2600
rect 14792 -2668 14856 -2634
rect 14792 -2702 14818 -2668
rect 14852 -2702 14856 -2668
rect 14792 -2736 14856 -2702
rect 14792 -2770 14818 -2736
rect 14852 -2770 14856 -2736
rect 14792 -2804 14856 -2770
rect 14792 -2838 14818 -2804
rect 14852 -2838 14856 -2804
rect 14792 -2872 14856 -2838
rect 14792 -2906 14818 -2872
rect 14852 -2906 14856 -2872
rect 14792 -2960 14856 -2906
<< psubdiffcont >>
rect 12598 -3524 12632 -3490
rect 12598 -3592 12632 -3558
rect 12598 -3660 12632 -3626
rect 12598 -3728 12632 -3694
rect 12598 -3796 12632 -3762
rect 12598 -3864 12632 -3830
rect 12598 -3932 12632 -3898
rect 12598 -4000 12632 -3966
rect 12598 -4068 12632 -4034
rect 12598 -4136 12632 -4102
rect 12598 -4204 12632 -4170
rect 12598 -4272 12632 -4238
rect 12598 -4340 12632 -4306
rect 12598 -4408 12632 -4374
rect 12934 -3498 12968 -3464
rect 12934 -3566 12968 -3532
rect 12934 -3634 12968 -3600
rect 12934 -3702 12968 -3668
rect 12934 -3770 12968 -3736
rect 12934 -3838 12968 -3804
rect 12934 -3906 12968 -3872
rect 12934 -3974 12968 -3940
rect 12934 -4042 12968 -4008
rect 12934 -4110 12968 -4076
rect 12934 -4178 12968 -4144
rect 12934 -4246 12968 -4212
rect 12934 -4314 12968 -4280
rect 12934 -4382 12968 -4348
rect 13270 -3498 13304 -3464
rect 13270 -3566 13304 -3532
rect 13270 -3634 13304 -3600
rect 13270 -3702 13304 -3668
rect 13270 -3770 13304 -3736
rect 13270 -3838 13304 -3804
rect 13270 -3906 13304 -3872
rect 13270 -3974 13304 -3940
rect 13270 -4042 13304 -4008
rect 13270 -4110 13304 -4076
rect 13270 -4178 13304 -4144
rect 13270 -4246 13304 -4212
rect 13270 -4314 13304 -4280
rect 13270 -4382 13304 -4348
rect 13606 -3498 13640 -3464
rect 13606 -3566 13640 -3532
rect 13606 -3634 13640 -3600
rect 13606 -3702 13640 -3668
rect 13606 -3770 13640 -3736
rect 13606 -3838 13640 -3804
rect 13606 -3906 13640 -3872
rect 13606 -3974 13640 -3940
rect 13606 -4042 13640 -4008
rect 13606 -4110 13640 -4076
rect 13606 -4178 13640 -4144
rect 13606 -4246 13640 -4212
rect 13606 -4314 13640 -4280
rect 13606 -4382 13640 -4348
rect 13942 -3498 13976 -3464
rect 13942 -3566 13976 -3532
rect 13942 -3634 13976 -3600
rect 13942 -3702 13976 -3668
rect 13942 -3770 13976 -3736
rect 13942 -3838 13976 -3804
rect 13942 -3906 13976 -3872
rect 13942 -3974 13976 -3940
rect 13942 -4042 13976 -4008
rect 13942 -4110 13976 -4076
rect 13942 -4178 13976 -4144
rect 13942 -4246 13976 -4212
rect 13942 -4314 13976 -4280
rect 13942 -4382 13976 -4348
rect 14278 -3498 14312 -3464
rect 14278 -3566 14312 -3532
rect 14278 -3634 14312 -3600
rect 14278 -3702 14312 -3668
rect 14278 -3770 14312 -3736
rect 14278 -3838 14312 -3804
rect 14278 -3906 14312 -3872
rect 14278 -3974 14312 -3940
rect 14278 -4042 14312 -4008
rect 14278 -4110 14312 -4076
rect 14278 -4178 14312 -4144
rect 14278 -4246 14312 -4212
rect 14278 -4314 14312 -4280
rect 14278 -4382 14312 -4348
rect 14614 -3498 14648 -3464
rect 14614 -3566 14648 -3532
rect 14614 -3634 14648 -3600
rect 14614 -3702 14648 -3668
rect 14614 -3770 14648 -3736
rect 14614 -3838 14648 -3804
rect 14614 -3906 14648 -3872
rect 14614 -3974 14648 -3940
rect 14614 -4042 14648 -4008
rect 14614 -4110 14648 -4076
rect 14614 -4178 14648 -4144
rect 14614 -4246 14648 -4212
rect 14614 -4314 14648 -4280
rect 14614 -4382 14648 -4348
<< nsubdiffcont >>
rect 12394 -2048 12428 -2014
rect 12394 -2116 12428 -2082
rect 12394 -2184 12428 -2150
rect 12394 -2252 12428 -2218
rect 12394 -2320 12428 -2286
rect 12394 -2388 12428 -2354
rect 12394 -2456 12428 -2422
rect 12394 -2524 12428 -2490
rect 12394 -2592 12428 -2558
rect 12394 -2660 12428 -2626
rect 12394 -2728 12428 -2694
rect 12394 -2796 12428 -2762
rect 12394 -2864 12428 -2830
rect 12394 -2932 12428 -2898
rect 12798 -2022 12832 -1988
rect 12798 -2090 12832 -2056
rect 12798 -2158 12832 -2124
rect 12798 -2226 12832 -2192
rect 12798 -2294 12832 -2260
rect 12798 -2362 12832 -2328
rect 12798 -2430 12832 -2396
rect 12798 -2498 12832 -2464
rect 12798 -2566 12832 -2532
rect 12798 -2634 12832 -2600
rect 12798 -2702 12832 -2668
rect 12798 -2770 12832 -2736
rect 12798 -2838 12832 -2804
rect 12798 -2906 12832 -2872
rect 13202 -2022 13236 -1988
rect 13202 -2090 13236 -2056
rect 13202 -2158 13236 -2124
rect 13202 -2226 13236 -2192
rect 13202 -2294 13236 -2260
rect 13202 -2362 13236 -2328
rect 13202 -2430 13236 -2396
rect 13202 -2498 13236 -2464
rect 13202 -2566 13236 -2532
rect 13202 -2634 13236 -2600
rect 13202 -2702 13236 -2668
rect 13202 -2770 13236 -2736
rect 13202 -2838 13236 -2804
rect 13202 -2906 13236 -2872
rect 13606 -2022 13640 -1988
rect 13606 -2090 13640 -2056
rect 13606 -2158 13640 -2124
rect 13606 -2226 13640 -2192
rect 13606 -2294 13640 -2260
rect 13606 -2362 13640 -2328
rect 13606 -2430 13640 -2396
rect 13606 -2498 13640 -2464
rect 13606 -2566 13640 -2532
rect 13606 -2634 13640 -2600
rect 13606 -2702 13640 -2668
rect 13606 -2770 13640 -2736
rect 13606 -2838 13640 -2804
rect 13606 -2906 13640 -2872
rect 14010 -2022 14044 -1988
rect 14010 -2090 14044 -2056
rect 14010 -2158 14044 -2124
rect 14010 -2226 14044 -2192
rect 14010 -2294 14044 -2260
rect 14010 -2362 14044 -2328
rect 14010 -2430 14044 -2396
rect 14010 -2498 14044 -2464
rect 14010 -2566 14044 -2532
rect 14010 -2634 14044 -2600
rect 14010 -2702 14044 -2668
rect 14010 -2770 14044 -2736
rect 14010 -2838 14044 -2804
rect 14010 -2906 14044 -2872
rect 14414 -2022 14448 -1988
rect 14414 -2090 14448 -2056
rect 14414 -2158 14448 -2124
rect 14414 -2226 14448 -2192
rect 14414 -2294 14448 -2260
rect 14414 -2362 14448 -2328
rect 14414 -2430 14448 -2396
rect 14414 -2498 14448 -2464
rect 14414 -2566 14448 -2532
rect 14414 -2634 14448 -2600
rect 14414 -2702 14448 -2668
rect 14414 -2770 14448 -2736
rect 14414 -2838 14448 -2804
rect 14414 -2906 14448 -2872
rect 14818 -2022 14852 -1988
rect 14818 -2090 14852 -2056
rect 14818 -2158 14852 -2124
rect 14818 -2226 14852 -2192
rect 14818 -2294 14852 -2260
rect 14818 -2362 14852 -2328
rect 14818 -2430 14852 -2396
rect 14818 -2498 14852 -2464
rect 14818 -2566 14852 -2532
rect 14818 -2634 14852 -2600
rect 14818 -2702 14852 -2668
rect 14818 -2770 14852 -2736
rect 14818 -2838 14852 -2804
rect 14818 -2906 14852 -2872
<< poly >>
rect 12768 -3414 12798 -3348
rect 13104 -3414 13134 -3348
rect 13440 -3414 13470 -3348
rect 13776 -3414 13806 -3348
rect 14112 -3414 14142 -3348
rect 14448 -3414 14478 -3348
rect 12768 -4524 12798 -4458
rect 13104 -4524 13134 -4458
rect 13440 -4524 13470 -4458
rect 13776 -4524 13806 -4458
rect 14112 -4524 14142 -4458
rect 14448 -4524 14478 -4458
<< locali >>
rect 12394 -1972 12428 -1956
rect 12394 -2964 12428 -2948
rect 12798 -1972 12832 -1956
rect 12798 -2964 12832 -2948
rect 13202 -1972 13236 -1956
rect 13202 -2964 13236 -2948
rect 13606 -1972 13640 -1956
rect 13606 -2964 13640 -2948
rect 14010 -1972 14044 -1956
rect 14010 -2964 14044 -2948
rect 14414 -1972 14448 -1956
rect 14414 -2964 14448 -2948
rect 14818 -1972 14852 -1956
rect 14818 -2964 14852 -2948
rect 12768 -3398 12798 -3364
rect 13104 -3398 13134 -3364
rect 13440 -3398 13470 -3364
rect 13776 -3398 13806 -3364
rect 14112 -3398 14142 -3364
rect 14448 -3398 14478 -3364
rect 12598 -3448 12632 -3432
rect 12598 -4440 12632 -4424
rect 12934 -3448 12968 -3432
rect 12934 -4440 12968 -4424
rect 13270 -3448 13304 -3432
rect 13270 -4440 13304 -4424
rect 13606 -3448 13640 -3432
rect 13606 -4440 13640 -4424
rect 13942 -3448 13976 -3432
rect 13942 -4440 13976 -4424
rect 14278 -3448 14312 -3432
rect 14278 -4440 14312 -4424
rect 14614 -3448 14648 -3432
rect 14614 -4440 14648 -4424
rect 12768 -4508 12798 -4474
rect 13104 -4508 13134 -4474
rect 13440 -4508 13470 -4474
rect 13776 -4508 13806 -4474
rect 14112 -4508 14142 -4474
rect 14448 -4508 14478 -4474
<< viali >>
rect 12394 -2014 12428 -1972
rect 12394 -2048 12428 -2014
rect 12394 -2082 12428 -2048
rect 12394 -2116 12428 -2082
rect 12394 -2150 12428 -2116
rect 12394 -2184 12428 -2150
rect 12394 -2218 12428 -2184
rect 12394 -2252 12428 -2218
rect 12394 -2286 12428 -2252
rect 12394 -2320 12428 -2286
rect 12394 -2354 12428 -2320
rect 12394 -2388 12428 -2354
rect 12394 -2422 12428 -2388
rect 12394 -2456 12428 -2422
rect 12394 -2490 12428 -2456
rect 12394 -2524 12428 -2490
rect 12394 -2558 12428 -2524
rect 12394 -2592 12428 -2558
rect 12394 -2626 12428 -2592
rect 12394 -2660 12428 -2626
rect 12394 -2694 12428 -2660
rect 12394 -2728 12428 -2694
rect 12394 -2762 12428 -2728
rect 12394 -2796 12428 -2762
rect 12394 -2830 12428 -2796
rect 12394 -2864 12428 -2830
rect 12394 -2898 12428 -2864
rect 12394 -2932 12428 -2898
rect 12394 -2948 12428 -2932
rect 12798 -1988 12832 -1972
rect 12798 -2022 12832 -1988
rect 12798 -2056 12832 -2022
rect 12798 -2090 12832 -2056
rect 12798 -2124 12832 -2090
rect 12798 -2158 12832 -2124
rect 12798 -2192 12832 -2158
rect 12798 -2226 12832 -2192
rect 12798 -2260 12832 -2226
rect 12798 -2294 12832 -2260
rect 12798 -2328 12832 -2294
rect 12798 -2362 12832 -2328
rect 12798 -2396 12832 -2362
rect 12798 -2430 12832 -2396
rect 12798 -2464 12832 -2430
rect 12798 -2498 12832 -2464
rect 12798 -2532 12832 -2498
rect 12798 -2566 12832 -2532
rect 12798 -2600 12832 -2566
rect 12798 -2634 12832 -2600
rect 12798 -2668 12832 -2634
rect 12798 -2702 12832 -2668
rect 12798 -2736 12832 -2702
rect 12798 -2770 12832 -2736
rect 12798 -2804 12832 -2770
rect 12798 -2838 12832 -2804
rect 12798 -2872 12832 -2838
rect 12798 -2906 12832 -2872
rect 12798 -2948 12832 -2906
rect 13202 -1988 13236 -1972
rect 13202 -2022 13236 -1988
rect 13202 -2056 13236 -2022
rect 13202 -2090 13236 -2056
rect 13202 -2124 13236 -2090
rect 13202 -2158 13236 -2124
rect 13202 -2192 13236 -2158
rect 13202 -2226 13236 -2192
rect 13202 -2260 13236 -2226
rect 13202 -2294 13236 -2260
rect 13202 -2328 13236 -2294
rect 13202 -2362 13236 -2328
rect 13202 -2396 13236 -2362
rect 13202 -2430 13236 -2396
rect 13202 -2464 13236 -2430
rect 13202 -2498 13236 -2464
rect 13202 -2532 13236 -2498
rect 13202 -2566 13236 -2532
rect 13202 -2600 13236 -2566
rect 13202 -2634 13236 -2600
rect 13202 -2668 13236 -2634
rect 13202 -2702 13236 -2668
rect 13202 -2736 13236 -2702
rect 13202 -2770 13236 -2736
rect 13202 -2804 13236 -2770
rect 13202 -2838 13236 -2804
rect 13202 -2872 13236 -2838
rect 13202 -2906 13236 -2872
rect 13202 -2948 13236 -2906
rect 13606 -1988 13640 -1972
rect 13606 -2022 13640 -1988
rect 13606 -2056 13640 -2022
rect 13606 -2090 13640 -2056
rect 13606 -2124 13640 -2090
rect 13606 -2158 13640 -2124
rect 13606 -2192 13640 -2158
rect 13606 -2226 13640 -2192
rect 13606 -2260 13640 -2226
rect 13606 -2294 13640 -2260
rect 13606 -2328 13640 -2294
rect 13606 -2362 13640 -2328
rect 13606 -2396 13640 -2362
rect 13606 -2430 13640 -2396
rect 13606 -2464 13640 -2430
rect 13606 -2498 13640 -2464
rect 13606 -2532 13640 -2498
rect 13606 -2566 13640 -2532
rect 13606 -2600 13640 -2566
rect 13606 -2634 13640 -2600
rect 13606 -2668 13640 -2634
rect 13606 -2702 13640 -2668
rect 13606 -2736 13640 -2702
rect 13606 -2770 13640 -2736
rect 13606 -2804 13640 -2770
rect 13606 -2838 13640 -2804
rect 13606 -2872 13640 -2838
rect 13606 -2906 13640 -2872
rect 13606 -2948 13640 -2906
rect 14010 -1988 14044 -1972
rect 14010 -2022 14044 -1988
rect 14010 -2056 14044 -2022
rect 14010 -2090 14044 -2056
rect 14010 -2124 14044 -2090
rect 14010 -2158 14044 -2124
rect 14010 -2192 14044 -2158
rect 14010 -2226 14044 -2192
rect 14010 -2260 14044 -2226
rect 14010 -2294 14044 -2260
rect 14010 -2328 14044 -2294
rect 14010 -2362 14044 -2328
rect 14010 -2396 14044 -2362
rect 14010 -2430 14044 -2396
rect 14010 -2464 14044 -2430
rect 14010 -2498 14044 -2464
rect 14010 -2532 14044 -2498
rect 14010 -2566 14044 -2532
rect 14010 -2600 14044 -2566
rect 14010 -2634 14044 -2600
rect 14010 -2668 14044 -2634
rect 14010 -2702 14044 -2668
rect 14010 -2736 14044 -2702
rect 14010 -2770 14044 -2736
rect 14010 -2804 14044 -2770
rect 14010 -2838 14044 -2804
rect 14010 -2872 14044 -2838
rect 14010 -2906 14044 -2872
rect 14010 -2948 14044 -2906
rect 14414 -1988 14448 -1972
rect 14414 -2022 14448 -1988
rect 14414 -2056 14448 -2022
rect 14414 -2090 14448 -2056
rect 14414 -2124 14448 -2090
rect 14414 -2158 14448 -2124
rect 14414 -2192 14448 -2158
rect 14414 -2226 14448 -2192
rect 14414 -2260 14448 -2226
rect 14414 -2294 14448 -2260
rect 14414 -2328 14448 -2294
rect 14414 -2362 14448 -2328
rect 14414 -2396 14448 -2362
rect 14414 -2430 14448 -2396
rect 14414 -2464 14448 -2430
rect 14414 -2498 14448 -2464
rect 14414 -2532 14448 -2498
rect 14414 -2566 14448 -2532
rect 14414 -2600 14448 -2566
rect 14414 -2634 14448 -2600
rect 14414 -2668 14448 -2634
rect 14414 -2702 14448 -2668
rect 14414 -2736 14448 -2702
rect 14414 -2770 14448 -2736
rect 14414 -2804 14448 -2770
rect 14414 -2838 14448 -2804
rect 14414 -2872 14448 -2838
rect 14414 -2906 14448 -2872
rect 14414 -2948 14448 -2906
rect 14818 -1988 14852 -1972
rect 14818 -2022 14852 -1988
rect 14818 -2056 14852 -2022
rect 14818 -2090 14852 -2056
rect 14818 -2124 14852 -2090
rect 14818 -2158 14852 -2124
rect 14818 -2192 14852 -2158
rect 14818 -2226 14852 -2192
rect 14818 -2260 14852 -2226
rect 14818 -2294 14852 -2260
rect 14818 -2328 14852 -2294
rect 14818 -2362 14852 -2328
rect 14818 -2396 14852 -2362
rect 14818 -2430 14852 -2396
rect 14818 -2464 14852 -2430
rect 14818 -2498 14852 -2464
rect 14818 -2532 14852 -2498
rect 14818 -2566 14852 -2532
rect 14818 -2600 14852 -2566
rect 14818 -2634 14852 -2600
rect 14818 -2668 14852 -2634
rect 14818 -2702 14852 -2668
rect 14818 -2736 14852 -2702
rect 14818 -2770 14852 -2736
rect 14818 -2804 14852 -2770
rect 14818 -2838 14852 -2804
rect 14818 -2872 14852 -2838
rect 14818 -2906 14852 -2872
rect 14818 -2948 14852 -2906
rect 12598 -3490 12632 -3448
rect 12598 -3524 12632 -3490
rect 12598 -3558 12632 -3524
rect 12598 -3592 12632 -3558
rect 12598 -3626 12632 -3592
rect 12598 -3660 12632 -3626
rect 12598 -3694 12632 -3660
rect 12598 -3728 12632 -3694
rect 12598 -3762 12632 -3728
rect 12598 -3796 12632 -3762
rect 12598 -3830 12632 -3796
rect 12598 -3864 12632 -3830
rect 12598 -3898 12632 -3864
rect 12598 -3932 12632 -3898
rect 12598 -3966 12632 -3932
rect 12598 -4000 12632 -3966
rect 12598 -4034 12632 -4000
rect 12598 -4068 12632 -4034
rect 12598 -4102 12632 -4068
rect 12598 -4136 12632 -4102
rect 12598 -4170 12632 -4136
rect 12598 -4204 12632 -4170
rect 12598 -4238 12632 -4204
rect 12598 -4272 12632 -4238
rect 12598 -4306 12632 -4272
rect 12598 -4340 12632 -4306
rect 12598 -4374 12632 -4340
rect 12598 -4408 12632 -4374
rect 12598 -4424 12632 -4408
rect 12934 -3464 12968 -3448
rect 12934 -3498 12968 -3464
rect 12934 -3532 12968 -3498
rect 12934 -3566 12968 -3532
rect 12934 -3600 12968 -3566
rect 12934 -3634 12968 -3600
rect 12934 -3668 12968 -3634
rect 12934 -3702 12968 -3668
rect 12934 -3736 12968 -3702
rect 12934 -3770 12968 -3736
rect 12934 -3804 12968 -3770
rect 12934 -3838 12968 -3804
rect 12934 -3872 12968 -3838
rect 12934 -3906 12968 -3872
rect 12934 -3940 12968 -3906
rect 12934 -3974 12968 -3940
rect 12934 -4008 12968 -3974
rect 12934 -4042 12968 -4008
rect 12934 -4076 12968 -4042
rect 12934 -4110 12968 -4076
rect 12934 -4144 12968 -4110
rect 12934 -4178 12968 -4144
rect 12934 -4212 12968 -4178
rect 12934 -4246 12968 -4212
rect 12934 -4280 12968 -4246
rect 12934 -4314 12968 -4280
rect 12934 -4348 12968 -4314
rect 12934 -4382 12968 -4348
rect 12934 -4424 12968 -4382
rect 13270 -3464 13304 -3448
rect 13270 -3498 13304 -3464
rect 13270 -3532 13304 -3498
rect 13270 -3566 13304 -3532
rect 13270 -3600 13304 -3566
rect 13270 -3634 13304 -3600
rect 13270 -3668 13304 -3634
rect 13270 -3702 13304 -3668
rect 13270 -3736 13304 -3702
rect 13270 -3770 13304 -3736
rect 13270 -3804 13304 -3770
rect 13270 -3838 13304 -3804
rect 13270 -3872 13304 -3838
rect 13270 -3906 13304 -3872
rect 13270 -3940 13304 -3906
rect 13270 -3974 13304 -3940
rect 13270 -4008 13304 -3974
rect 13270 -4042 13304 -4008
rect 13270 -4076 13304 -4042
rect 13270 -4110 13304 -4076
rect 13270 -4144 13304 -4110
rect 13270 -4178 13304 -4144
rect 13270 -4212 13304 -4178
rect 13270 -4246 13304 -4212
rect 13270 -4280 13304 -4246
rect 13270 -4314 13304 -4280
rect 13270 -4348 13304 -4314
rect 13270 -4382 13304 -4348
rect 13270 -4424 13304 -4382
rect 13606 -3464 13640 -3448
rect 13606 -3498 13640 -3464
rect 13606 -3532 13640 -3498
rect 13606 -3566 13640 -3532
rect 13606 -3600 13640 -3566
rect 13606 -3634 13640 -3600
rect 13606 -3668 13640 -3634
rect 13606 -3702 13640 -3668
rect 13606 -3736 13640 -3702
rect 13606 -3770 13640 -3736
rect 13606 -3804 13640 -3770
rect 13606 -3838 13640 -3804
rect 13606 -3872 13640 -3838
rect 13606 -3906 13640 -3872
rect 13606 -3940 13640 -3906
rect 13606 -3974 13640 -3940
rect 13606 -4008 13640 -3974
rect 13606 -4042 13640 -4008
rect 13606 -4076 13640 -4042
rect 13606 -4110 13640 -4076
rect 13606 -4144 13640 -4110
rect 13606 -4178 13640 -4144
rect 13606 -4212 13640 -4178
rect 13606 -4246 13640 -4212
rect 13606 -4280 13640 -4246
rect 13606 -4314 13640 -4280
rect 13606 -4348 13640 -4314
rect 13606 -4382 13640 -4348
rect 13606 -4424 13640 -4382
rect 13942 -3464 13976 -3448
rect 13942 -3498 13976 -3464
rect 13942 -3532 13976 -3498
rect 13942 -3566 13976 -3532
rect 13942 -3600 13976 -3566
rect 13942 -3634 13976 -3600
rect 13942 -3668 13976 -3634
rect 13942 -3702 13976 -3668
rect 13942 -3736 13976 -3702
rect 13942 -3770 13976 -3736
rect 13942 -3804 13976 -3770
rect 13942 -3838 13976 -3804
rect 13942 -3872 13976 -3838
rect 13942 -3906 13976 -3872
rect 13942 -3940 13976 -3906
rect 13942 -3974 13976 -3940
rect 13942 -4008 13976 -3974
rect 13942 -4042 13976 -4008
rect 13942 -4076 13976 -4042
rect 13942 -4110 13976 -4076
rect 13942 -4144 13976 -4110
rect 13942 -4178 13976 -4144
rect 13942 -4212 13976 -4178
rect 13942 -4246 13976 -4212
rect 13942 -4280 13976 -4246
rect 13942 -4314 13976 -4280
rect 13942 -4348 13976 -4314
rect 13942 -4382 13976 -4348
rect 13942 -4424 13976 -4382
rect 14278 -3464 14312 -3448
rect 14278 -3498 14312 -3464
rect 14278 -3532 14312 -3498
rect 14278 -3566 14312 -3532
rect 14278 -3600 14312 -3566
rect 14278 -3634 14312 -3600
rect 14278 -3668 14312 -3634
rect 14278 -3702 14312 -3668
rect 14278 -3736 14312 -3702
rect 14278 -3770 14312 -3736
rect 14278 -3804 14312 -3770
rect 14278 -3838 14312 -3804
rect 14278 -3872 14312 -3838
rect 14278 -3906 14312 -3872
rect 14278 -3940 14312 -3906
rect 14278 -3974 14312 -3940
rect 14278 -4008 14312 -3974
rect 14278 -4042 14312 -4008
rect 14278 -4076 14312 -4042
rect 14278 -4110 14312 -4076
rect 14278 -4144 14312 -4110
rect 14278 -4178 14312 -4144
rect 14278 -4212 14312 -4178
rect 14278 -4246 14312 -4212
rect 14278 -4280 14312 -4246
rect 14278 -4314 14312 -4280
rect 14278 -4348 14312 -4314
rect 14278 -4382 14312 -4348
rect 14278 -4424 14312 -4382
rect 14614 -3464 14648 -3448
rect 14614 -3498 14648 -3464
rect 14614 -3532 14648 -3498
rect 14614 -3566 14648 -3532
rect 14614 -3600 14648 -3566
rect 14614 -3634 14648 -3600
rect 14614 -3668 14648 -3634
rect 14614 -3702 14648 -3668
rect 14614 -3736 14648 -3702
rect 14614 -3770 14648 -3736
rect 14614 -3804 14648 -3770
rect 14614 -3838 14648 -3804
rect 14614 -3872 14648 -3838
rect 14614 -3906 14648 -3872
rect 14614 -3940 14648 -3906
rect 14614 -3974 14648 -3940
rect 14614 -4008 14648 -3974
rect 14614 -4042 14648 -4008
rect 14614 -4076 14648 -4042
rect 14614 -4110 14648 -4076
rect 14614 -4144 14648 -4110
rect 14614 -4178 14648 -4144
rect 14614 -4212 14648 -4178
rect 14614 -4246 14648 -4212
rect 14614 -4280 14648 -4246
rect 14614 -4314 14648 -4280
rect 14614 -4348 14648 -4314
rect 14614 -4382 14648 -4348
rect 14614 -4424 14648 -4382
<< metal1 >>
rect 12234 -1498 12346 -1488
rect 12234 -1666 12264 -1498
rect 12320 -1666 12346 -1498
rect 11974 -4558 12198 -1798
rect 12234 -3248 12346 -1666
rect 12374 -1768 15182 -1762
rect 12374 -1820 12394 -1768
rect 15174 -1820 15182 -1768
rect 12374 -1826 15182 -1820
rect 12374 -1972 12486 -1826
rect 12516 -1920 12710 -1872
rect 12374 -2948 12394 -1972
rect 12428 -2948 12486 -1972
rect 12374 -2960 12486 -2948
rect 12584 -1972 12642 -1962
rect 12584 -2954 12642 -2948
rect 12758 -1972 12870 -1826
rect 12920 -1920 13114 -1872
rect 12758 -2948 12798 -1972
rect 12832 -2948 12870 -1972
rect 12758 -2960 12870 -2948
rect 12988 -1972 13046 -1962
rect 12988 -2954 13046 -2948
rect 13162 -1972 13274 -1826
rect 13324 -1920 13518 -1872
rect 13162 -2948 13202 -1972
rect 13236 -2948 13274 -1972
rect 13162 -2960 13274 -2948
rect 13392 -1972 13450 -1962
rect 13392 -2954 13450 -2948
rect 13566 -1972 13678 -1826
rect 13728 -1920 13922 -1872
rect 13566 -2948 13606 -1972
rect 13640 -2948 13678 -1972
rect 13566 -2960 13678 -2948
rect 13796 -1972 13854 -1962
rect 13796 -2954 13854 -2948
rect 13970 -1972 14082 -1826
rect 14132 -1920 14326 -1872
rect 13970 -2948 14010 -1972
rect 14044 -2948 14082 -1972
rect 13970 -2960 14082 -2948
rect 14200 -1972 14258 -1962
rect 14200 -2954 14258 -2948
rect 14374 -1972 14486 -1826
rect 14536 -1920 14730 -1872
rect 14374 -2948 14414 -1972
rect 14448 -2948 14486 -1972
rect 14374 -2960 14486 -2948
rect 14604 -1972 14662 -1962
rect 14604 -2954 14662 -2948
rect 14758 -1972 14870 -1826
rect 14758 -2948 14818 -1972
rect 14852 -2948 14870 -1972
rect 14758 -2960 14870 -2948
rect 12516 -3060 12710 -3000
rect 12920 -3060 13114 -3000
rect 12588 -3102 12710 -3060
rect 12588 -3108 12838 -3102
rect 12812 -3160 12838 -3108
rect 12588 -3166 12838 -3160
rect 12234 -3306 12346 -3300
rect 12704 -3348 12838 -3166
rect 12950 -3242 13084 -3060
rect 13324 -3102 13518 -3000
rect 13324 -3108 13548 -3102
rect 13324 -3166 13548 -3160
rect 12950 -3248 13198 -3242
rect 13174 -3300 13198 -3248
rect 12950 -3306 13198 -3300
rect 12704 -3404 12862 -3348
rect 13040 -3404 13198 -3306
rect 13376 -3404 13534 -3166
rect 13728 -3242 13922 -3000
rect 14132 -3102 14326 -3000
rect 14078 -3108 14326 -3102
rect 14302 -3160 14326 -3108
rect 14078 -3166 14326 -3160
rect 14536 -3078 14730 -3000
rect 13704 -3248 13928 -3242
rect 13704 -3306 13928 -3300
rect 13712 -3404 13870 -3306
rect 14078 -3348 14190 -3166
rect 14536 -3242 14656 -3078
rect 14424 -3248 14656 -3242
rect 14648 -3300 14656 -3248
rect 14424 -3306 14656 -3300
rect 14764 -3108 14876 -3102
rect 14424 -3348 14542 -3306
rect 14048 -3404 14206 -3348
rect 14384 -3404 14542 -3348
rect 12560 -3448 12672 -3436
rect 12560 -4424 12598 -3448
rect 12632 -4424 12672 -3448
rect 12560 -4558 12672 -4424
rect 12754 -3446 12812 -3434
rect 12754 -4436 12812 -4422
rect 12894 -3448 13006 -3436
rect 12894 -4424 12934 -3448
rect 12968 -4424 13006 -3448
rect 12704 -4514 12862 -4468
rect 12894 -4558 13006 -4424
rect 13090 -3446 13148 -3434
rect 13090 -4436 13148 -4422
rect 13230 -3448 13342 -3436
rect 13230 -4424 13270 -3448
rect 13304 -4424 13342 -3448
rect 13040 -4514 13198 -4468
rect 13230 -4558 13342 -4424
rect 13426 -3446 13484 -3434
rect 13426 -4436 13484 -4422
rect 13566 -3448 13678 -3436
rect 13566 -4424 13606 -3448
rect 13640 -4424 13678 -3448
rect 13376 -4514 13534 -4468
rect 13566 -4558 13678 -4424
rect 13762 -3446 13820 -3434
rect 13762 -4436 13820 -4422
rect 13902 -3448 14014 -3436
rect 13902 -4424 13942 -3448
rect 13976 -4424 14014 -3448
rect 13712 -4514 13870 -4468
rect 13902 -4558 14014 -4424
rect 14098 -3446 14156 -3434
rect 14098 -4436 14156 -4422
rect 14238 -3448 14350 -3436
rect 14238 -4424 14278 -3448
rect 14312 -4424 14350 -3448
rect 14048 -4514 14206 -4468
rect 14238 -4558 14350 -4424
rect 14434 -3446 14492 -3434
rect 14434 -4436 14492 -4422
rect 14572 -3448 14684 -3434
rect 14572 -4424 14614 -3448
rect 14648 -4424 14684 -3448
rect 14384 -4514 14542 -4468
rect 14572 -4558 14684 -4424
rect 11974 -4564 14684 -4558
rect 11974 -4616 11982 -4564
rect 14664 -4616 14684 -4564
rect 11974 -4622 14684 -4616
rect 11974 -4646 12198 -4622
rect 14764 -4708 14876 -3160
rect 14958 -4668 15182 -1826
rect 14764 -4876 14792 -4708
rect 14848 -4876 14876 -4708
rect 14764 -4886 14876 -4876
<< via1 >>
rect 12264 -1666 12320 -1498
rect 12394 -1820 15174 -1768
rect 12584 -2948 12642 -1972
rect 12988 -2948 13046 -1972
rect 13392 -2948 13450 -1972
rect 13796 -2948 13854 -1972
rect 14200 -2948 14258 -1972
rect 14604 -2948 14662 -1972
rect 12588 -3160 12812 -3108
rect 12234 -3300 12346 -3248
rect 13324 -3160 13548 -3108
rect 12950 -3300 13174 -3248
rect 14078 -3160 14302 -3108
rect 13704 -3300 13928 -3248
rect 14424 -3300 14648 -3248
rect 14764 -3160 14876 -3108
rect 12754 -4422 12812 -3446
rect 13090 -4422 13148 -3446
rect 13426 -4422 13484 -3446
rect 13762 -4422 13820 -3446
rect 14098 -4422 14156 -3446
rect 14434 -4422 14492 -3446
rect 11982 -4616 14664 -4564
rect 14792 -4876 14848 -4708
<< metal2 >>
rect 12234 -1498 12346 -1488
rect 12234 -1666 12264 -1498
rect 12320 -1666 12346 -1498
rect 12234 -1676 12346 -1666
rect 12374 -1768 15182 -1738
rect 12374 -1820 12394 -1768
rect 15174 -1820 15182 -1768
rect 12374 -1850 15182 -1820
rect 12584 -1972 12642 -1962
rect 12584 -2960 12642 -2948
rect 12988 -1972 13046 -1962
rect 12988 -2960 13046 -2948
rect 13392 -1972 13450 -1962
rect 13392 -2960 13450 -2948
rect 13796 -1972 13854 -1962
rect 13796 -2960 13854 -2948
rect 14200 -1972 14258 -1962
rect 14200 -2960 14258 -2948
rect 14604 -1972 14662 -1962
rect 14604 -2960 14662 -2948
rect 12588 -3078 12710 -3050
rect 12510 -3108 14876 -3078
rect 12510 -3160 12588 -3108
rect 12812 -3160 13324 -3108
rect 13548 -3160 14078 -3108
rect 14302 -3160 14764 -3108
rect 12510 -3190 14876 -3160
rect 12234 -3248 14736 -3218
rect 12346 -3300 12950 -3248
rect 13174 -3300 13704 -3248
rect 13928 -3300 14424 -3248
rect 14648 -3300 14736 -3248
rect 12234 -3330 14736 -3300
rect 12754 -3446 12812 -3434
rect 12754 -4436 12812 -4422
rect 13090 -3446 13148 -3434
rect 13090 -4436 13148 -4422
rect 13426 -3446 13484 -3434
rect 13426 -4436 13484 -4422
rect 13762 -3446 13820 -3434
rect 13762 -4436 13820 -4422
rect 14098 -3446 14156 -3434
rect 14098 -4436 14156 -4422
rect 14434 -3446 14492 -3434
rect 14434 -4436 14492 -4422
rect 11974 -4564 14684 -4534
rect 11974 -4616 11982 -4564
rect 14664 -4616 14684 -4564
rect 11974 -4646 14684 -4616
rect 14764 -4708 14876 -4698
rect 14764 -4876 14792 -4708
rect 14848 -4876 14876 -4708
rect 14764 -4886 14876 -4876
<< via2 >>
rect 12264 -1666 12320 -1498
rect 12584 -2948 12642 -1972
rect 12988 -2948 13046 -1972
rect 13392 -2948 13450 -1972
rect 13796 -2948 13854 -1972
rect 14200 -2948 14258 -1972
rect 14604 -2948 14662 -1972
rect 12754 -4422 12812 -3446
rect 13090 -4422 13148 -3446
rect 13426 -4422 13484 -3446
rect 13762 -4422 13820 -3446
rect 14098 -4422 14156 -3446
rect 14434 -4422 14492 -3446
rect 14792 -4876 14848 -4708
<< metal3 >>
rect 11974 -1498 15182 -1464
rect 11974 -1544 12264 -1498
rect 12320 -1544 15182 -1498
rect 11974 -1614 11980 -1544
rect 15176 -1614 15182 -1544
rect 11974 -1666 12264 -1614
rect 12320 -1666 15182 -1614
rect 11974 -1694 15182 -1666
rect 12578 -1972 12758 -1694
rect 12578 -2948 12584 -1972
rect 12642 -2948 12758 -1972
rect 12578 -3440 12758 -2948
rect 12982 -1972 13162 -1960
rect 12982 -2948 12988 -1972
rect 13046 -2948 13162 -1972
rect 12578 -3446 12818 -3440
rect 12578 -4422 12754 -3446
rect 12812 -4422 12818 -3446
rect 12578 -4428 12818 -4422
rect 12982 -3446 13162 -2948
rect 12982 -4422 13090 -3446
rect 13148 -4422 13162 -3446
rect 12982 -4682 13162 -4422
rect 13386 -1972 13566 -1694
rect 13386 -2948 13392 -1972
rect 13450 -2948 13566 -1972
rect 13386 -3446 13566 -2948
rect 13386 -4422 13426 -3446
rect 13484 -4422 13566 -3446
rect 13386 -4428 13566 -4422
rect 13740 -1972 13920 -1960
rect 13740 -2948 13796 -1972
rect 13854 -2948 13920 -1972
rect 13740 -3446 13920 -2948
rect 13740 -4422 13762 -3446
rect 13820 -4422 13920 -3446
rect 13740 -4682 13920 -4422
rect 14084 -1972 14264 -1694
rect 14084 -2948 14200 -1972
rect 14258 -2948 14264 -1972
rect 14084 -3446 14264 -2948
rect 14084 -4422 14098 -3446
rect 14156 -4422 14264 -3446
rect 14084 -4428 14264 -4422
rect 14428 -1972 14668 -1960
rect 14428 -2948 14604 -1972
rect 14662 -2948 14668 -1972
rect 14428 -2960 14668 -2948
rect 14428 -3446 14614 -2960
rect 14428 -4422 14434 -3446
rect 14492 -4422 14614 -3446
rect 14428 -4682 14614 -4422
rect 11974 -4708 15182 -4682
rect 11974 -4766 14792 -4708
rect 14848 -4766 15182 -4708
rect 11974 -4836 11980 -4766
rect 15176 -4836 15182 -4766
rect 11974 -4876 14792 -4836
rect 14848 -4876 15182 -4836
rect 11974 -11464 15182 -4876
<< via3 >>
rect 11980 -1614 12264 -1544
rect 12264 -1614 12320 -1544
rect 12320 -1614 15176 -1544
rect 11980 -4836 14792 -4766
rect 14792 -4836 14848 -4766
rect 14848 -4836 15176 -4766
<< metal4 >>
rect 11974 -1544 15182 5906
rect 11974 -1614 11980 -1544
rect 15176 -1614 15182 -1544
rect 11974 -1620 15182 -1614
rect 11974 -4766 15182 -4760
rect 11974 -4836 11980 -4766
rect 15176 -4836 15182 -4766
rect 11974 -12424 15182 -4836
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M11
timestamp 1680265380
transform -1 0 12736 0 1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M12
timestamp 1680265380
transform 1 0 12830 0 -1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M13
timestamp 1680265380
transform -1 0 13408 0 1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M14
timestamp 1680265380
transform 1 0 13502 0 -1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M15
timestamp 1680265380
transform -1 0 14080 0 1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M16
timestamp 1680265380
transform 1 0 14174 0 -1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M21
timestamp 1680265380
transform -1 0 13072 0 1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M22
timestamp 1680265380
transform 1 0 13166 0 -1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M23
timestamp 1680265380
transform -1 0 13744 0 1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M24
timestamp 1680265380
transform 1 0 13838 0 -1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M25
timestamp 1680265380
transform -1 0 14416 0 1 -3936
box -76 -588 76 588
use sky130_fd_pr__nfet_01v8_lvt_R7Y3EQ  M26
timestamp 1680265380
transform 1 0 14510 0 -1 -3936
box -76 -588 76 588
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M31
timestamp 1680265380
transform -1 0 12549 0 1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M32
timestamp 1680265380
transform 1 0 12677 0 -1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M33
timestamp 1680265380
transform -1 0 13357 0 1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M34
timestamp 1680265380
transform 1 0 13485 0 -1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M35
timestamp 1680265380
transform -1 0 14165 0 1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M36
timestamp 1680265380
transform 1 0 14293 0 -1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M41
timestamp 1680265380
transform -1 0 12953 0 1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M42
timestamp 1680265380
transform 1 0 13081 0 -1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M43
timestamp 1680265380
transform -1 0 13761 0 1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M44
timestamp 1680265380
transform 1 0 13889 0 -1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M45
timestamp 1680265380
transform -1 0 14569 0 1 -2460
box -129 -600 129 600
use sky130_fd_pr__pfet_01v8_lvt_4QFV24  M46
timestamp 1680265380
transform 1 0 14697 0 -1 -2460
box -129 -600 129 600
<< labels >>
flabel metal1 14958 -4668 15182 -1864 0 FreeMono 1280 90 0 0 out2
port 3 nsew
flabel metal1 11974 -4514 12198 -1798 0 FreeMono 1280 90 0 0 vss
port 2 nsew
flabel metal4 11974 -12424 15182 -11464 0 FreeMono 1600 0 0 0 vinn
port 1 nsew
flabel metal4 11974 4946 15182 5906 0 FreeMono 1600 0 0 0 vinp
port 0 nsew
<< end >>
