magic
tech sky130A
magscale 1 2
timestamp 1680213737
<< pwell >>
rect -201 -668 201 668
<< psubdiff >>
rect -165 598 -69 632
rect 69 598 165 632
rect -165 536 -131 598
rect 131 536 165 598
rect -165 -598 -131 -536
rect 131 -598 165 -536
rect -165 -632 -69 -598
rect 69 -632 165 -598
<< psubdiffcont >>
rect -69 598 69 632
rect -165 -536 -131 536
rect 131 -536 165 536
rect -69 -632 69 -598
<< xpolycontact >>
rect -35 70 35 502
rect -35 -502 35 -70
<< xpolyres >>
rect -35 -70 35 70
<< locali >>
rect -165 598 -69 632
rect 69 598 165 632
rect -165 536 -131 598
rect 131 536 165 598
rect -165 -598 -131 -536
rect 131 -598 165 -536
rect -165 -632 -69 -598
rect 69 -632 165 -598
<< viali >>
rect -19 87 19 484
rect -19 -484 19 -87
<< metal1 >>
rect -25 484 25 496
rect -25 87 -19 484
rect 19 87 25 484
rect -25 75 25 87
rect -25 -87 25 -75
rect -25 -484 -19 -87
rect 19 -484 25 -87
rect -25 -496 25 -484
<< res0p35 >>
rect -37 -72 37 72
<< properties >>
string FIXED_BBOX -148 -615 148 615
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.350 l 0.7 m 1 nx 1 wmin 0.350 lmin 0.50 rho 2000 val 5.075k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
