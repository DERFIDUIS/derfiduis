magic
tech sky130A
magscale 1 2
timestamp 1681575212
<< nwell >>
rect 1894 86 1960 212
rect 3518 86 3584 212
rect 5140 170 5206 212
rect 5140 112 5276 170
rect 5140 86 5206 112
rect 1894 52 1968 86
rect 3518 52 3592 86
rect 5140 52 5214 86
rect 1894 18 1960 52
rect 3518 18 3584 52
rect 5140 18 5206 52
rect 1894 -16 1968 18
rect 3518 -16 3592 18
rect 5140 -16 5214 18
rect 1894 -50 1960 -16
rect 3518 -50 3584 -16
rect 5140 -50 5206 -16
rect 1894 -84 1968 -50
rect 3518 -84 3592 -50
rect 5140 -84 5214 -50
rect 1894 -118 1960 -84
rect 3518 -118 3584 -84
rect 5140 -118 5206 -84
rect 1894 -152 1968 -118
rect 3518 -152 3592 -118
rect 5140 -152 5214 -118
rect 1894 -186 1960 -152
rect 3518 -186 3584 -152
rect 5140 -186 5206 -152
rect 1894 -220 1968 -186
rect 3518 -220 3592 -186
rect 5140 -220 5214 -186
rect 1894 -254 1960 -220
rect 3518 -254 3584 -220
rect 5140 -254 5206 -220
rect 1894 -288 1968 -254
rect 3518 -288 3592 -254
rect 5140 -288 5214 -254
rect 1894 -322 1960 -288
rect 3518 -322 3584 -288
rect 5140 -322 5206 -288
rect 1894 -356 1968 -322
rect 3518 -356 3592 -322
rect 5140 -356 5214 -322
rect 1894 -390 1960 -356
rect 3518 -390 3584 -356
rect 5140 -390 5206 -356
rect 1894 -424 1968 -390
rect 3518 -424 3592 -390
rect 5140 -424 5214 -390
rect 1894 -458 1960 -424
rect 3518 -458 3584 -424
rect 5140 -458 5206 -424
rect 1894 -492 1968 -458
rect 3518 -492 3592 -458
rect 5140 -492 5214 -458
rect 1894 -526 1960 -492
rect 3518 -526 3584 -492
rect 5140 -526 5206 -492
rect 1894 -560 1968 -526
rect 3518 -560 3592 -526
rect 5140 -560 5214 -526
rect 1894 -594 1960 -560
rect 3518 -594 3584 -560
rect 5140 -594 5206 -560
rect 1894 -628 1968 -594
rect 3518 -628 3592 -594
rect 5140 -628 5214 -594
rect 1894 -662 1960 -628
rect 3518 -662 3584 -628
rect 5140 -662 5206 -628
rect 1894 -696 1968 -662
rect 3518 -696 3592 -662
rect 5140 -696 5214 -662
rect 1894 -730 1960 -696
rect 3518 -730 3584 -696
rect 5140 -730 5206 -696
rect 1894 -764 1968 -730
rect 3518 -764 3592 -730
rect 5140 -764 5214 -730
rect 1894 -798 1960 -764
rect 3518 -798 3584 -764
rect 5140 -798 5206 -764
rect 1894 -832 1968 -798
rect 3518 -832 3592 -798
rect 5140 -832 5214 -798
rect 1894 -866 1960 -832
rect 3518 -866 3584 -832
rect 5140 -866 5206 -832
rect 1894 -900 1968 -866
rect 3518 -900 3592 -866
rect 5140 -900 5214 -866
rect 1894 -934 1960 -900
rect 3518 -934 3584 -900
rect 5140 -934 5206 -900
rect 1894 -968 1968 -934
rect 3518 -968 3592 -934
rect 5140 -968 5214 -934
rect 1894 -1002 1960 -968
rect 3518 -1002 3584 -968
rect 5140 -1002 5206 -968
rect 1894 -1036 1968 -1002
rect 3518 -1036 3592 -1002
rect 5140 -1036 5214 -1002
rect 1894 -1070 1960 -1036
rect 3518 -1070 3584 -1036
rect 5140 -1070 5206 -1036
rect 1894 -1104 1968 -1070
rect 3518 -1104 3592 -1070
rect 5140 -1104 5214 -1070
rect 1894 -1138 1960 -1104
rect 3518 -1138 3584 -1104
rect 5140 -1138 5206 -1104
rect 1894 -1172 1968 -1138
rect 3518 -1172 3592 -1138
rect 5140 -1172 5214 -1138
rect 1894 -1206 1960 -1172
rect 3518 -1206 3584 -1172
rect 5140 -1206 5206 -1172
rect 1894 -1240 1968 -1206
rect 3518 -1240 3592 -1206
rect 5140 -1240 5214 -1206
rect 1894 -1274 1960 -1240
rect 3518 -1274 3584 -1240
rect 5140 -1274 5206 -1240
rect 1894 -1308 1968 -1274
rect 3518 -1308 3592 -1274
rect 5140 -1308 5214 -1274
rect 1894 -1342 1960 -1308
rect 3518 -1342 3584 -1308
rect 5140 -1342 5206 -1308
rect 1894 -1376 1968 -1342
rect 3518 -1376 3592 -1342
rect 5140 -1376 5214 -1342
rect 1894 -1410 1960 -1376
rect 3518 -1410 3584 -1376
rect 5140 -1410 5206 -1376
rect 1894 -1444 1968 -1410
rect 3518 -1444 3592 -1410
rect 5140 -1444 5214 -1410
rect 1894 -1478 1960 -1444
rect 3518 -1478 3584 -1444
rect 5140 -1478 5206 -1444
rect 1894 -1512 1968 -1478
rect 3518 -1512 3592 -1478
rect 5140 -1512 5214 -1478
rect 1894 -1546 1960 -1512
rect 3518 -1546 3584 -1512
rect 5140 -1546 5206 -1512
rect 1894 -1580 1968 -1546
rect 3518 -1580 3592 -1546
rect 5140 -1580 5214 -1546
rect 1894 -1614 1960 -1580
rect 3518 -1614 3584 -1580
rect 5140 -1614 5206 -1580
rect 1894 -1648 1968 -1614
rect 3518 -1648 3592 -1614
rect 5140 -1648 5214 -1614
rect 1894 -1682 1960 -1648
rect 3518 -1682 3584 -1648
rect 5140 -1682 5206 -1648
rect 1894 -1716 1968 -1682
rect 3518 -1716 3592 -1682
rect 5140 -1716 5214 -1682
rect 1894 -1750 1960 -1716
rect 3518 -1750 3584 -1716
rect 5140 -1750 5206 -1716
rect 1894 -1784 1968 -1750
rect 3518 -1784 3592 -1750
rect 5140 -1784 5214 -1750
rect 1894 -1818 1960 -1784
rect 3518 -1818 3584 -1784
rect 5140 -1818 5206 -1784
rect 1894 -1852 1968 -1818
rect 3518 -1852 3592 -1818
rect 5140 -1852 5214 -1818
rect 1894 -1886 1960 -1852
rect 3518 -1886 3584 -1852
rect 5140 -1886 5206 -1852
rect 1894 -1920 1968 -1886
rect 3518 -1920 3592 -1886
rect 5140 -1920 5214 -1886
rect 1894 -1954 1960 -1920
rect 3518 -1954 3584 -1920
rect 5140 -1954 5206 -1920
rect 1894 -1988 1968 -1954
rect 3518 -1988 3592 -1954
rect 5140 -1988 5214 -1954
rect 1894 -2022 1960 -1988
rect 3518 -2022 3584 -1988
rect 5140 -2022 5206 -1988
rect 1894 -2056 1968 -2022
rect 3518 -2056 3592 -2022
rect 5140 -2056 5214 -2022
rect 1894 -2090 1960 -2056
rect 3518 -2090 3584 -2056
rect 5140 -2090 5206 -2056
rect 1894 -2124 1968 -2090
rect 3518 -2124 3592 -2090
rect 5140 -2124 5214 -2090
rect 1894 -2158 1960 -2124
rect 3518 -2158 3584 -2124
rect 5140 -2158 5206 -2124
rect 1894 -2192 1968 -2158
rect 3518 -2192 3592 -2158
rect 5140 -2192 5214 -2158
rect 1894 -2388 1960 -2192
rect 3518 -2388 3584 -2192
rect 5140 -2388 5206 -2192
rect 2007 -3443 3273 -3416
rect 3611 -3443 4877 -3413
rect 5232 -3443 6498 -3413
rect 2007 -4652 3273 -4625
rect 3611 -4655 4877 -4625
rect 5232 -4655 6498 -4625
<< ndiff >>
rect 1994 -3316 1996 -2516
rect 3618 -3316 3620 -2516
rect 5240 -3316 5242 -2516
<< pdiff >>
rect 1994 -2288 1996 112
rect 3618 -2288 3620 112
rect 5240 -2288 5242 112
<< psubdiff >>
rect 1930 -2574 1994 -2516
rect 1930 -2608 1934 -2574
rect 1968 -2608 1994 -2574
rect 1930 -2642 1994 -2608
rect 1930 -2676 1934 -2642
rect 1968 -2676 1994 -2642
rect 1930 -2710 1994 -2676
rect 1930 -2744 1934 -2710
rect 1968 -2744 1994 -2710
rect 1930 -2778 1994 -2744
rect 1930 -2812 1934 -2778
rect 1968 -2812 1994 -2778
rect 1930 -2846 1994 -2812
rect 1930 -2880 1934 -2846
rect 1968 -2880 1994 -2846
rect 1930 -2914 1994 -2880
rect 1930 -2948 1934 -2914
rect 1968 -2948 1994 -2914
rect 1930 -2982 1994 -2948
rect 1930 -3016 1934 -2982
rect 1968 -3016 1994 -2982
rect 1930 -3050 1994 -3016
rect 1930 -3084 1934 -3050
rect 1968 -3084 1994 -3050
rect 1930 -3118 1994 -3084
rect 1930 -3152 1934 -3118
rect 1968 -3152 1994 -3118
rect 1930 -3186 1994 -3152
rect 1930 -3220 1934 -3186
rect 1968 -3220 1994 -3186
rect 1930 -3254 1994 -3220
rect 1930 -3288 1934 -3254
rect 1968 -3288 1994 -3254
rect 1930 -3316 1994 -3288
rect 3554 -2574 3618 -2516
rect 3554 -2608 3558 -2574
rect 3592 -2608 3618 -2574
rect 3554 -2642 3618 -2608
rect 3554 -2676 3558 -2642
rect 3592 -2676 3618 -2642
rect 3554 -2710 3618 -2676
rect 3554 -2744 3558 -2710
rect 3592 -2744 3618 -2710
rect 3554 -2778 3618 -2744
rect 3554 -2812 3558 -2778
rect 3592 -2812 3618 -2778
rect 3554 -2846 3618 -2812
rect 3554 -2880 3558 -2846
rect 3592 -2880 3618 -2846
rect 3554 -2914 3618 -2880
rect 3554 -2948 3558 -2914
rect 3592 -2948 3618 -2914
rect 3554 -2982 3618 -2948
rect 3554 -3016 3558 -2982
rect 3592 -3016 3618 -2982
rect 3554 -3050 3618 -3016
rect 3554 -3084 3558 -3050
rect 3592 -3084 3618 -3050
rect 3554 -3118 3618 -3084
rect 3554 -3152 3558 -3118
rect 3592 -3152 3618 -3118
rect 3554 -3186 3618 -3152
rect 3554 -3220 3558 -3186
rect 3592 -3220 3618 -3186
rect 3554 -3254 3618 -3220
rect 3554 -3288 3558 -3254
rect 3592 -3288 3618 -3254
rect 3554 -3316 3618 -3288
rect 5176 -2574 5240 -2516
rect 5176 -2608 5180 -2574
rect 5214 -2608 5240 -2574
rect 5176 -2642 5240 -2608
rect 5176 -2676 5180 -2642
rect 5214 -2676 5240 -2642
rect 5176 -2710 5240 -2676
rect 5176 -2744 5180 -2710
rect 5214 -2744 5240 -2710
rect 5176 -2778 5240 -2744
rect 5176 -2812 5180 -2778
rect 5214 -2812 5240 -2778
rect 5176 -2846 5240 -2812
rect 5176 -2880 5180 -2846
rect 5214 -2880 5240 -2846
rect 5176 -2914 5240 -2880
rect 5176 -2948 5180 -2914
rect 5214 -2948 5240 -2914
rect 5176 -2982 5240 -2948
rect 5176 -3016 5180 -2982
rect 5214 -3016 5240 -2982
rect 5176 -3050 5240 -3016
rect 5176 -3084 5180 -3050
rect 5214 -3084 5240 -3050
rect 5176 -3118 5240 -3084
rect 5176 -3152 5180 -3118
rect 5214 -3152 5240 -3118
rect 5176 -3186 5240 -3152
rect 5176 -3220 5180 -3186
rect 5214 -3220 5240 -3186
rect 5176 -3254 5240 -3220
rect 5176 -3288 5180 -3254
rect 5214 -3288 5240 -3254
rect 5176 -3316 5240 -3288
rect 1925 -3592 1981 -3534
rect 1925 -3626 1933 -3592
rect 1967 -3626 1981 -3592
rect 1925 -3660 1981 -3626
rect 1925 -3694 1933 -3660
rect 1967 -3694 1981 -3660
rect 1925 -3728 1981 -3694
rect 1925 -3762 1933 -3728
rect 1967 -3762 1981 -3728
rect 1925 -3796 1981 -3762
rect 1925 -3830 1933 -3796
rect 1967 -3830 1981 -3796
rect 1925 -3864 1981 -3830
rect 1925 -3898 1933 -3864
rect 1967 -3898 1981 -3864
rect 1925 -3932 1981 -3898
rect 1925 -3966 1933 -3932
rect 1967 -3966 1981 -3932
rect 1925 -4000 1981 -3966
rect 1925 -4034 1933 -4000
rect 1967 -4034 1981 -4000
rect 1925 -4068 1981 -4034
rect 1925 -4102 1933 -4068
rect 1967 -4102 1981 -4068
rect 1925 -4136 1981 -4102
rect 1925 -4170 1933 -4136
rect 1967 -4170 1981 -4136
rect 1925 -4204 1981 -4170
rect 1925 -4238 1933 -4204
rect 1967 -4238 1981 -4204
rect 1925 -4272 1981 -4238
rect 1925 -4306 1933 -4272
rect 1967 -4306 1981 -4272
rect 1925 -4340 1981 -4306
rect 1925 -4374 1933 -4340
rect 1967 -4374 1981 -4340
rect 1925 -4408 1981 -4374
rect 1925 -4442 1933 -4408
rect 1967 -4442 1981 -4408
rect 1925 -4476 1981 -4442
rect 1925 -4510 1933 -4476
rect 1967 -4510 1981 -4476
rect 1925 -4534 1981 -4510
rect 3527 -3592 3583 -3534
rect 3527 -3626 3535 -3592
rect 3569 -3626 3583 -3592
rect 3527 -3660 3583 -3626
rect 3527 -3694 3535 -3660
rect 3569 -3694 3583 -3660
rect 3527 -3728 3583 -3694
rect 3527 -3762 3535 -3728
rect 3569 -3762 3583 -3728
rect 3527 -3796 3583 -3762
rect 3527 -3830 3535 -3796
rect 3569 -3830 3583 -3796
rect 3527 -3864 3583 -3830
rect 3527 -3898 3535 -3864
rect 3569 -3898 3583 -3864
rect 3527 -3932 3583 -3898
rect 3527 -3966 3535 -3932
rect 3569 -3966 3583 -3932
rect 3527 -4000 3583 -3966
rect 3527 -4034 3535 -4000
rect 3569 -4034 3583 -4000
rect 3527 -4068 3583 -4034
rect 3527 -4102 3535 -4068
rect 3569 -4102 3583 -4068
rect 3527 -4136 3583 -4102
rect 3527 -4170 3535 -4136
rect 3569 -4170 3583 -4136
rect 3527 -4204 3583 -4170
rect 3527 -4238 3535 -4204
rect 3569 -4238 3583 -4204
rect 3527 -4272 3583 -4238
rect 3527 -4306 3535 -4272
rect 3569 -4306 3583 -4272
rect 3527 -4340 3583 -4306
rect 3527 -4374 3535 -4340
rect 3569 -4374 3583 -4340
rect 3527 -4408 3583 -4374
rect 3527 -4442 3535 -4408
rect 3569 -4442 3583 -4408
rect 3527 -4476 3583 -4442
rect 3527 -4510 3535 -4476
rect 3569 -4510 3583 -4476
rect 3527 -4534 3583 -4510
rect 5150 -3592 5206 -3534
rect 5150 -3626 5158 -3592
rect 5192 -3626 5206 -3592
rect 5150 -3660 5206 -3626
rect 5150 -3694 5158 -3660
rect 5192 -3694 5206 -3660
rect 5150 -3728 5206 -3694
rect 5150 -3762 5158 -3728
rect 5192 -3762 5206 -3728
rect 5150 -3796 5206 -3762
rect 5150 -3830 5158 -3796
rect 5192 -3830 5206 -3796
rect 5150 -3864 5206 -3830
rect 5150 -3898 5158 -3864
rect 5192 -3898 5206 -3864
rect 5150 -3932 5206 -3898
rect 5150 -3966 5158 -3932
rect 5192 -3966 5206 -3932
rect 5150 -4000 5206 -3966
rect 5150 -4034 5158 -4000
rect 5192 -4034 5206 -4000
rect 5150 -4068 5206 -4034
rect 5150 -4102 5158 -4068
rect 5192 -4102 5206 -4068
rect 5150 -4136 5206 -4102
rect 5150 -4170 5158 -4136
rect 5192 -4170 5206 -4136
rect 5150 -4204 5206 -4170
rect 5150 -4238 5158 -4204
rect 5192 -4238 5206 -4204
rect 5150 -4272 5206 -4238
rect 5150 -4306 5158 -4272
rect 5192 -4306 5206 -4272
rect 5150 -4340 5206 -4306
rect 5150 -4374 5158 -4340
rect 5192 -4374 5206 -4340
rect 5150 -4408 5206 -4374
rect 5150 -4442 5158 -4408
rect 5192 -4442 5206 -4408
rect 5150 -4476 5206 -4442
rect 5150 -4510 5158 -4476
rect 5192 -4510 5206 -4476
rect 5150 -4534 5206 -4510
<< nsubdiff >>
rect 1930 86 1994 112
rect 1930 52 1934 86
rect 1968 52 1994 86
rect 1930 18 1994 52
rect 1930 -16 1934 18
rect 1968 -16 1994 18
rect 1930 -50 1994 -16
rect 1930 -84 1934 -50
rect 1968 -84 1994 -50
rect 1930 -118 1994 -84
rect 1930 -152 1934 -118
rect 1968 -152 1994 -118
rect 1930 -186 1994 -152
rect 1930 -220 1934 -186
rect 1968 -220 1994 -186
rect 1930 -254 1994 -220
rect 1930 -288 1934 -254
rect 1968 -288 1994 -254
rect 1930 -322 1994 -288
rect 1930 -356 1934 -322
rect 1968 -356 1994 -322
rect 1930 -390 1994 -356
rect 1930 -424 1934 -390
rect 1968 -424 1994 -390
rect 1930 -458 1994 -424
rect 1930 -492 1934 -458
rect 1968 -492 1994 -458
rect 1930 -526 1994 -492
rect 1930 -560 1934 -526
rect 1968 -560 1994 -526
rect 1930 -594 1994 -560
rect 1930 -628 1934 -594
rect 1968 -628 1994 -594
rect 1930 -662 1994 -628
rect 1930 -696 1934 -662
rect 1968 -696 1994 -662
rect 1930 -730 1994 -696
rect 1930 -764 1934 -730
rect 1968 -764 1994 -730
rect 1930 -798 1994 -764
rect 1930 -832 1934 -798
rect 1968 -832 1994 -798
rect 1930 -866 1994 -832
rect 1930 -900 1934 -866
rect 1968 -900 1994 -866
rect 1930 -934 1994 -900
rect 1930 -968 1934 -934
rect 1968 -968 1994 -934
rect 1930 -1002 1994 -968
rect 1930 -1036 1934 -1002
rect 1968 -1036 1994 -1002
rect 1930 -1070 1994 -1036
rect 1930 -1104 1934 -1070
rect 1968 -1104 1994 -1070
rect 1930 -1138 1994 -1104
rect 1930 -1172 1934 -1138
rect 1968 -1172 1994 -1138
rect 1930 -1206 1994 -1172
rect 1930 -1240 1934 -1206
rect 1968 -1240 1994 -1206
rect 1930 -1274 1994 -1240
rect 1930 -1308 1934 -1274
rect 1968 -1308 1994 -1274
rect 1930 -1342 1994 -1308
rect 1930 -1376 1934 -1342
rect 1968 -1376 1994 -1342
rect 1930 -1410 1994 -1376
rect 1930 -1444 1934 -1410
rect 1968 -1444 1994 -1410
rect 1930 -1478 1994 -1444
rect 1930 -1512 1934 -1478
rect 1968 -1512 1994 -1478
rect 1930 -1546 1994 -1512
rect 1930 -1580 1934 -1546
rect 1968 -1580 1994 -1546
rect 1930 -1614 1994 -1580
rect 1930 -1648 1934 -1614
rect 1968 -1648 1994 -1614
rect 1930 -1682 1994 -1648
rect 1930 -1716 1934 -1682
rect 1968 -1716 1994 -1682
rect 1930 -1750 1994 -1716
rect 1930 -1784 1934 -1750
rect 1968 -1784 1994 -1750
rect 1930 -1818 1994 -1784
rect 1930 -1852 1934 -1818
rect 1968 -1852 1994 -1818
rect 1930 -1886 1994 -1852
rect 1930 -1920 1934 -1886
rect 1968 -1920 1994 -1886
rect 1930 -1954 1994 -1920
rect 1930 -1988 1934 -1954
rect 1968 -1988 1994 -1954
rect 1930 -2022 1994 -1988
rect 1930 -2056 1934 -2022
rect 1968 -2056 1994 -2022
rect 1930 -2090 1994 -2056
rect 1930 -2124 1934 -2090
rect 1968 -2124 1994 -2090
rect 1930 -2158 1994 -2124
rect 1930 -2192 1934 -2158
rect 1968 -2192 1994 -2158
rect 1930 -2226 1994 -2192
rect 1930 -2260 1934 -2226
rect 1968 -2260 1994 -2226
rect 1930 -2288 1994 -2260
rect 3554 86 3618 112
rect 3554 52 3558 86
rect 3592 52 3618 86
rect 3554 18 3618 52
rect 3554 -16 3558 18
rect 3592 -16 3618 18
rect 3554 -50 3618 -16
rect 3554 -84 3558 -50
rect 3592 -84 3618 -50
rect 3554 -118 3618 -84
rect 3554 -152 3558 -118
rect 3592 -152 3618 -118
rect 3554 -186 3618 -152
rect 3554 -220 3558 -186
rect 3592 -220 3618 -186
rect 3554 -254 3618 -220
rect 3554 -288 3558 -254
rect 3592 -288 3618 -254
rect 3554 -322 3618 -288
rect 3554 -356 3558 -322
rect 3592 -356 3618 -322
rect 3554 -390 3618 -356
rect 3554 -424 3558 -390
rect 3592 -424 3618 -390
rect 3554 -458 3618 -424
rect 3554 -492 3558 -458
rect 3592 -492 3618 -458
rect 3554 -526 3618 -492
rect 3554 -560 3558 -526
rect 3592 -560 3618 -526
rect 3554 -594 3618 -560
rect 3554 -628 3558 -594
rect 3592 -628 3618 -594
rect 3554 -662 3618 -628
rect 3554 -696 3558 -662
rect 3592 -696 3618 -662
rect 3554 -730 3618 -696
rect 3554 -764 3558 -730
rect 3592 -764 3618 -730
rect 3554 -798 3618 -764
rect 3554 -832 3558 -798
rect 3592 -832 3618 -798
rect 3554 -866 3618 -832
rect 3554 -900 3558 -866
rect 3592 -900 3618 -866
rect 3554 -934 3618 -900
rect 3554 -968 3558 -934
rect 3592 -968 3618 -934
rect 3554 -1002 3618 -968
rect 3554 -1036 3558 -1002
rect 3592 -1036 3618 -1002
rect 3554 -1070 3618 -1036
rect 3554 -1104 3558 -1070
rect 3592 -1104 3618 -1070
rect 3554 -1138 3618 -1104
rect 3554 -1172 3558 -1138
rect 3592 -1172 3618 -1138
rect 3554 -1206 3618 -1172
rect 3554 -1240 3558 -1206
rect 3592 -1240 3618 -1206
rect 3554 -1274 3618 -1240
rect 3554 -1308 3558 -1274
rect 3592 -1308 3618 -1274
rect 3554 -1342 3618 -1308
rect 3554 -1376 3558 -1342
rect 3592 -1376 3618 -1342
rect 3554 -1410 3618 -1376
rect 3554 -1444 3558 -1410
rect 3592 -1444 3618 -1410
rect 3554 -1478 3618 -1444
rect 3554 -1512 3558 -1478
rect 3592 -1512 3618 -1478
rect 3554 -1546 3618 -1512
rect 3554 -1580 3558 -1546
rect 3592 -1580 3618 -1546
rect 3554 -1614 3618 -1580
rect 3554 -1648 3558 -1614
rect 3592 -1648 3618 -1614
rect 3554 -1682 3618 -1648
rect 3554 -1716 3558 -1682
rect 3592 -1716 3618 -1682
rect 3554 -1750 3618 -1716
rect 3554 -1784 3558 -1750
rect 3592 -1784 3618 -1750
rect 3554 -1818 3618 -1784
rect 3554 -1852 3558 -1818
rect 3592 -1852 3618 -1818
rect 3554 -1886 3618 -1852
rect 3554 -1920 3558 -1886
rect 3592 -1920 3618 -1886
rect 3554 -1954 3618 -1920
rect 3554 -1988 3558 -1954
rect 3592 -1988 3618 -1954
rect 3554 -2022 3618 -1988
rect 3554 -2056 3558 -2022
rect 3592 -2056 3618 -2022
rect 3554 -2090 3618 -2056
rect 3554 -2124 3558 -2090
rect 3592 -2124 3618 -2090
rect 3554 -2158 3618 -2124
rect 3554 -2192 3558 -2158
rect 3592 -2192 3618 -2158
rect 3554 -2226 3618 -2192
rect 3554 -2260 3558 -2226
rect 3592 -2260 3618 -2226
rect 3554 -2288 3618 -2260
rect 5176 86 5240 112
rect 5176 52 5180 86
rect 5214 52 5240 86
rect 5176 18 5240 52
rect 5176 -16 5180 18
rect 5214 -16 5240 18
rect 5176 -50 5240 -16
rect 5176 -84 5180 -50
rect 5214 -84 5240 -50
rect 5176 -118 5240 -84
rect 5176 -152 5180 -118
rect 5214 -152 5240 -118
rect 5176 -186 5240 -152
rect 5176 -220 5180 -186
rect 5214 -220 5240 -186
rect 5176 -254 5240 -220
rect 5176 -288 5180 -254
rect 5214 -288 5240 -254
rect 5176 -322 5240 -288
rect 5176 -356 5180 -322
rect 5214 -356 5240 -322
rect 5176 -390 5240 -356
rect 5176 -424 5180 -390
rect 5214 -424 5240 -390
rect 5176 -458 5240 -424
rect 5176 -492 5180 -458
rect 5214 -492 5240 -458
rect 5176 -526 5240 -492
rect 5176 -560 5180 -526
rect 5214 -560 5240 -526
rect 5176 -594 5240 -560
rect 5176 -628 5180 -594
rect 5214 -628 5240 -594
rect 5176 -662 5240 -628
rect 5176 -696 5180 -662
rect 5214 -696 5240 -662
rect 5176 -730 5240 -696
rect 5176 -764 5180 -730
rect 5214 -764 5240 -730
rect 5176 -798 5240 -764
rect 5176 -832 5180 -798
rect 5214 -832 5240 -798
rect 5176 -866 5240 -832
rect 5176 -900 5180 -866
rect 5214 -900 5240 -866
rect 5176 -934 5240 -900
rect 5176 -968 5180 -934
rect 5214 -968 5240 -934
rect 5176 -1002 5240 -968
rect 5176 -1036 5180 -1002
rect 5214 -1036 5240 -1002
rect 5176 -1070 5240 -1036
rect 5176 -1104 5180 -1070
rect 5214 -1104 5240 -1070
rect 5176 -1138 5240 -1104
rect 5176 -1172 5180 -1138
rect 5214 -1172 5240 -1138
rect 5176 -1206 5240 -1172
rect 5176 -1240 5180 -1206
rect 5214 -1240 5240 -1206
rect 5176 -1274 5240 -1240
rect 5176 -1308 5180 -1274
rect 5214 -1308 5240 -1274
rect 5176 -1342 5240 -1308
rect 5176 -1376 5180 -1342
rect 5214 -1376 5240 -1342
rect 5176 -1410 5240 -1376
rect 5176 -1444 5180 -1410
rect 5214 -1444 5240 -1410
rect 5176 -1478 5240 -1444
rect 5176 -1512 5180 -1478
rect 5214 -1512 5240 -1478
rect 5176 -1546 5240 -1512
rect 5176 -1580 5180 -1546
rect 5214 -1580 5240 -1546
rect 5176 -1614 5240 -1580
rect 5176 -1648 5180 -1614
rect 5214 -1648 5240 -1614
rect 5176 -1682 5240 -1648
rect 5176 -1716 5180 -1682
rect 5214 -1716 5240 -1682
rect 5176 -1750 5240 -1716
rect 5176 -1784 5180 -1750
rect 5214 -1784 5240 -1750
rect 5176 -1818 5240 -1784
rect 5176 -1852 5180 -1818
rect 5214 -1852 5240 -1818
rect 5176 -1886 5240 -1852
rect 5176 -1920 5180 -1886
rect 5214 -1920 5240 -1886
rect 5176 -1954 5240 -1920
rect 5176 -1988 5180 -1954
rect 5214 -1988 5240 -1954
rect 5176 -2022 5240 -1988
rect 5176 -2056 5180 -2022
rect 5214 -2056 5240 -2022
rect 5176 -2090 5240 -2056
rect 5176 -2124 5180 -2090
rect 5214 -2124 5240 -2090
rect 5176 -2158 5240 -2124
rect 5176 -2192 5180 -2158
rect 5214 -2192 5240 -2158
rect 5176 -2226 5240 -2192
rect 5176 -2260 5180 -2226
rect 5214 -2260 5240 -2226
rect 5176 -2288 5240 -2260
<< psubdiffcont >>
rect 1934 -2608 1968 -2574
rect 1934 -2676 1968 -2642
rect 1934 -2744 1968 -2710
rect 1934 -2812 1968 -2778
rect 1934 -2880 1968 -2846
rect 1934 -2948 1968 -2914
rect 1934 -3016 1968 -2982
rect 1934 -3084 1968 -3050
rect 1934 -3152 1968 -3118
rect 1934 -3220 1968 -3186
rect 1934 -3288 1968 -3254
rect 3558 -2608 3592 -2574
rect 3558 -2676 3592 -2642
rect 3558 -2744 3592 -2710
rect 3558 -2812 3592 -2778
rect 3558 -2880 3592 -2846
rect 3558 -2948 3592 -2914
rect 3558 -3016 3592 -2982
rect 3558 -3084 3592 -3050
rect 3558 -3152 3592 -3118
rect 3558 -3220 3592 -3186
rect 3558 -3288 3592 -3254
rect 5180 -2608 5214 -2574
rect 5180 -2676 5214 -2642
rect 5180 -2744 5214 -2710
rect 5180 -2812 5214 -2778
rect 5180 -2880 5214 -2846
rect 5180 -2948 5214 -2914
rect 5180 -3016 5214 -2982
rect 5180 -3084 5214 -3050
rect 5180 -3152 5214 -3118
rect 5180 -3220 5214 -3186
rect 5180 -3288 5214 -3254
rect 1933 -3626 1967 -3592
rect 1933 -3694 1967 -3660
rect 1933 -3762 1967 -3728
rect 1933 -3830 1967 -3796
rect 1933 -3898 1967 -3864
rect 1933 -3966 1967 -3932
rect 1933 -4034 1967 -4000
rect 1933 -4102 1967 -4068
rect 1933 -4170 1967 -4136
rect 1933 -4238 1967 -4204
rect 1933 -4306 1967 -4272
rect 1933 -4374 1967 -4340
rect 1933 -4442 1967 -4408
rect 1933 -4510 1967 -4476
rect 3535 -3626 3569 -3592
rect 3535 -3694 3569 -3660
rect 3535 -3762 3569 -3728
rect 3535 -3830 3569 -3796
rect 3535 -3898 3569 -3864
rect 3535 -3966 3569 -3932
rect 3535 -4034 3569 -4000
rect 3535 -4102 3569 -4068
rect 3535 -4170 3569 -4136
rect 3535 -4238 3569 -4204
rect 3535 -4306 3569 -4272
rect 3535 -4374 3569 -4340
rect 3535 -4442 3569 -4408
rect 3535 -4510 3569 -4476
rect 5158 -3626 5192 -3592
rect 5158 -3694 5192 -3660
rect 5158 -3762 5192 -3728
rect 5158 -3830 5192 -3796
rect 5158 -3898 5192 -3864
rect 5158 -3966 5192 -3932
rect 5158 -4034 5192 -4000
rect 5158 -4102 5192 -4068
rect 5158 -4170 5192 -4136
rect 5158 -4238 5192 -4204
rect 5158 -4306 5192 -4272
rect 5158 -4374 5192 -4340
rect 5158 -4442 5192 -4408
rect 5158 -4510 5192 -4476
<< nsubdiffcont >>
rect 1934 52 1968 86
rect 1934 -16 1968 18
rect 1934 -84 1968 -50
rect 1934 -152 1968 -118
rect 1934 -220 1968 -186
rect 1934 -288 1968 -254
rect 1934 -356 1968 -322
rect 1934 -424 1968 -390
rect 1934 -492 1968 -458
rect 1934 -560 1968 -526
rect 1934 -628 1968 -594
rect 1934 -696 1968 -662
rect 1934 -764 1968 -730
rect 1934 -832 1968 -798
rect 1934 -900 1968 -866
rect 1934 -968 1968 -934
rect 1934 -1036 1968 -1002
rect 1934 -1104 1968 -1070
rect 1934 -1172 1968 -1138
rect 1934 -1240 1968 -1206
rect 1934 -1308 1968 -1274
rect 1934 -1376 1968 -1342
rect 1934 -1444 1968 -1410
rect 1934 -1512 1968 -1478
rect 1934 -1580 1968 -1546
rect 1934 -1648 1968 -1614
rect 1934 -1716 1968 -1682
rect 1934 -1784 1968 -1750
rect 1934 -1852 1968 -1818
rect 1934 -1920 1968 -1886
rect 1934 -1988 1968 -1954
rect 1934 -2056 1968 -2022
rect 1934 -2124 1968 -2090
rect 1934 -2192 1968 -2158
rect 1934 -2260 1968 -2226
rect 3558 52 3592 86
rect 3558 -16 3592 18
rect 3558 -84 3592 -50
rect 3558 -152 3592 -118
rect 3558 -220 3592 -186
rect 3558 -288 3592 -254
rect 3558 -356 3592 -322
rect 3558 -424 3592 -390
rect 3558 -492 3592 -458
rect 3558 -560 3592 -526
rect 3558 -628 3592 -594
rect 3558 -696 3592 -662
rect 3558 -764 3592 -730
rect 3558 -832 3592 -798
rect 3558 -900 3592 -866
rect 3558 -968 3592 -934
rect 3558 -1036 3592 -1002
rect 3558 -1104 3592 -1070
rect 3558 -1172 3592 -1138
rect 3558 -1240 3592 -1206
rect 3558 -1308 3592 -1274
rect 3558 -1376 3592 -1342
rect 3558 -1444 3592 -1410
rect 3558 -1512 3592 -1478
rect 3558 -1580 3592 -1546
rect 3558 -1648 3592 -1614
rect 3558 -1716 3592 -1682
rect 3558 -1784 3592 -1750
rect 3558 -1852 3592 -1818
rect 3558 -1920 3592 -1886
rect 3558 -1988 3592 -1954
rect 3558 -2056 3592 -2022
rect 3558 -2124 3592 -2090
rect 3558 -2192 3592 -2158
rect 3558 -2260 3592 -2226
rect 5180 52 5214 86
rect 5180 -16 5214 18
rect 5180 -84 5214 -50
rect 5180 -152 5214 -118
rect 5180 -220 5214 -186
rect 5180 -288 5214 -254
rect 5180 -356 5214 -322
rect 5180 -424 5214 -390
rect 5180 -492 5214 -458
rect 5180 -560 5214 -526
rect 5180 -628 5214 -594
rect 5180 -696 5214 -662
rect 5180 -764 5214 -730
rect 5180 -832 5214 -798
rect 5180 -900 5214 -866
rect 5180 -968 5214 -934
rect 5180 -1036 5214 -1002
rect 5180 -1104 5214 -1070
rect 5180 -1172 5214 -1138
rect 5180 -1240 5214 -1206
rect 5180 -1308 5214 -1274
rect 5180 -1376 5214 -1342
rect 5180 -1444 5214 -1410
rect 5180 -1512 5214 -1478
rect 5180 -1580 5214 -1546
rect 5180 -1648 5214 -1614
rect 5180 -1716 5214 -1682
rect 5180 -1784 5214 -1750
rect 5180 -1852 5214 -1818
rect 5180 -1920 5214 -1886
rect 5180 -1988 5214 -1954
rect 5180 -2056 5214 -2022
rect 5180 -2124 5214 -2090
rect 5180 -2192 5214 -2158
rect 5180 -2260 5214 -2226
<< locali >>
rect 1934 100 1968 116
rect 1934 -2292 1968 -2276
rect 3558 100 3592 116
rect 3558 -2292 3592 -2276
rect 5180 100 5214 116
rect 5180 -2292 5214 -2276
rect 1934 -2528 1968 -2512
rect 1934 -3320 1968 -3304
rect 3558 -2528 3592 -2512
rect 3558 -3320 3592 -3304
rect 5180 -2528 5214 -2512
rect 5180 -3320 5214 -3304
rect 1933 -3558 1967 -3542
rect 1933 -4526 1967 -4510
rect 3535 -3558 3569 -3542
rect 3535 -4526 3569 -4510
rect 5158 -3558 5192 -3542
rect 5158 -4526 5192 -4510
<< viali >>
rect 1934 86 1968 100
rect 1934 52 1968 86
rect 1934 18 1968 52
rect 1934 -16 1968 18
rect 1934 -50 1968 -16
rect 1934 -84 1968 -50
rect 1934 -118 1968 -84
rect 1934 -152 1968 -118
rect 1934 -186 1968 -152
rect 1934 -220 1968 -186
rect 1934 -254 1968 -220
rect 1934 -288 1968 -254
rect 1934 -322 1968 -288
rect 1934 -356 1968 -322
rect 1934 -390 1968 -356
rect 1934 -424 1968 -390
rect 1934 -458 1968 -424
rect 1934 -492 1968 -458
rect 1934 -526 1968 -492
rect 1934 -560 1968 -526
rect 1934 -594 1968 -560
rect 1934 -628 1968 -594
rect 1934 -662 1968 -628
rect 1934 -696 1968 -662
rect 1934 -730 1968 -696
rect 1934 -764 1968 -730
rect 1934 -798 1968 -764
rect 1934 -832 1968 -798
rect 1934 -866 1968 -832
rect 1934 -900 1968 -866
rect 1934 -934 1968 -900
rect 1934 -968 1968 -934
rect 1934 -1002 1968 -968
rect 1934 -1036 1968 -1002
rect 1934 -1070 1968 -1036
rect 1934 -1104 1968 -1070
rect 1934 -1138 1968 -1104
rect 1934 -1172 1968 -1138
rect 1934 -1206 1968 -1172
rect 1934 -1240 1968 -1206
rect 1934 -1274 1968 -1240
rect 1934 -1308 1968 -1274
rect 1934 -1342 1968 -1308
rect 1934 -1376 1968 -1342
rect 1934 -1410 1968 -1376
rect 1934 -1444 1968 -1410
rect 1934 -1478 1968 -1444
rect 1934 -1512 1968 -1478
rect 1934 -1546 1968 -1512
rect 1934 -1580 1968 -1546
rect 1934 -1614 1968 -1580
rect 1934 -1648 1968 -1614
rect 1934 -1682 1968 -1648
rect 1934 -1716 1968 -1682
rect 1934 -1750 1968 -1716
rect 1934 -1784 1968 -1750
rect 1934 -1818 1968 -1784
rect 1934 -1852 1968 -1818
rect 1934 -1886 1968 -1852
rect 1934 -1920 1968 -1886
rect 1934 -1954 1968 -1920
rect 1934 -1988 1968 -1954
rect 1934 -2022 1968 -1988
rect 1934 -2056 1968 -2022
rect 1934 -2090 1968 -2056
rect 1934 -2124 1968 -2090
rect 1934 -2158 1968 -2124
rect 1934 -2192 1968 -2158
rect 1934 -2226 1968 -2192
rect 1934 -2260 1968 -2226
rect 1934 -2276 1968 -2260
rect 3558 86 3592 100
rect 3558 52 3592 86
rect 3558 18 3592 52
rect 3558 -16 3592 18
rect 3558 -50 3592 -16
rect 3558 -84 3592 -50
rect 3558 -118 3592 -84
rect 3558 -152 3592 -118
rect 3558 -186 3592 -152
rect 3558 -220 3592 -186
rect 3558 -254 3592 -220
rect 3558 -288 3592 -254
rect 3558 -322 3592 -288
rect 3558 -356 3592 -322
rect 3558 -390 3592 -356
rect 3558 -424 3592 -390
rect 3558 -458 3592 -424
rect 3558 -492 3592 -458
rect 3558 -526 3592 -492
rect 3558 -560 3592 -526
rect 3558 -594 3592 -560
rect 3558 -628 3592 -594
rect 3558 -662 3592 -628
rect 3558 -696 3592 -662
rect 3558 -730 3592 -696
rect 3558 -764 3592 -730
rect 3558 -798 3592 -764
rect 3558 -832 3592 -798
rect 3558 -866 3592 -832
rect 3558 -900 3592 -866
rect 3558 -934 3592 -900
rect 3558 -968 3592 -934
rect 3558 -1002 3592 -968
rect 3558 -1036 3592 -1002
rect 3558 -1070 3592 -1036
rect 3558 -1104 3592 -1070
rect 3558 -1138 3592 -1104
rect 3558 -1172 3592 -1138
rect 3558 -1206 3592 -1172
rect 3558 -1240 3592 -1206
rect 3558 -1274 3592 -1240
rect 3558 -1308 3592 -1274
rect 3558 -1342 3592 -1308
rect 3558 -1376 3592 -1342
rect 3558 -1410 3592 -1376
rect 3558 -1444 3592 -1410
rect 3558 -1478 3592 -1444
rect 3558 -1512 3592 -1478
rect 3558 -1546 3592 -1512
rect 3558 -1580 3592 -1546
rect 3558 -1614 3592 -1580
rect 3558 -1648 3592 -1614
rect 3558 -1682 3592 -1648
rect 3558 -1716 3592 -1682
rect 3558 -1750 3592 -1716
rect 3558 -1784 3592 -1750
rect 3558 -1818 3592 -1784
rect 3558 -1852 3592 -1818
rect 3558 -1886 3592 -1852
rect 3558 -1920 3592 -1886
rect 3558 -1954 3592 -1920
rect 3558 -1988 3592 -1954
rect 3558 -2022 3592 -1988
rect 3558 -2056 3592 -2022
rect 3558 -2090 3592 -2056
rect 3558 -2124 3592 -2090
rect 3558 -2158 3592 -2124
rect 3558 -2192 3592 -2158
rect 3558 -2226 3592 -2192
rect 3558 -2260 3592 -2226
rect 3558 -2276 3592 -2260
rect 5180 86 5214 100
rect 5180 52 5214 86
rect 5180 18 5214 52
rect 5180 -16 5214 18
rect 5180 -50 5214 -16
rect 5180 -84 5214 -50
rect 5180 -118 5214 -84
rect 5180 -152 5214 -118
rect 5180 -186 5214 -152
rect 5180 -220 5214 -186
rect 5180 -254 5214 -220
rect 5180 -288 5214 -254
rect 5180 -322 5214 -288
rect 5180 -356 5214 -322
rect 5180 -390 5214 -356
rect 5180 -424 5214 -390
rect 5180 -458 5214 -424
rect 5180 -492 5214 -458
rect 5180 -526 5214 -492
rect 5180 -560 5214 -526
rect 5180 -594 5214 -560
rect 5180 -628 5214 -594
rect 5180 -662 5214 -628
rect 5180 -696 5214 -662
rect 5180 -730 5214 -696
rect 5180 -764 5214 -730
rect 5180 -798 5214 -764
rect 5180 -832 5214 -798
rect 5180 -866 5214 -832
rect 5180 -900 5214 -866
rect 5180 -934 5214 -900
rect 5180 -968 5214 -934
rect 5180 -1002 5214 -968
rect 5180 -1036 5214 -1002
rect 5180 -1070 5214 -1036
rect 5180 -1104 5214 -1070
rect 5180 -1138 5214 -1104
rect 5180 -1172 5214 -1138
rect 5180 -1206 5214 -1172
rect 5180 -1240 5214 -1206
rect 5180 -1274 5214 -1240
rect 5180 -1308 5214 -1274
rect 5180 -1342 5214 -1308
rect 5180 -1376 5214 -1342
rect 5180 -1410 5214 -1376
rect 5180 -1444 5214 -1410
rect 5180 -1478 5214 -1444
rect 5180 -1512 5214 -1478
rect 5180 -1546 5214 -1512
rect 5180 -1580 5214 -1546
rect 5180 -1614 5214 -1580
rect 5180 -1648 5214 -1614
rect 5180 -1682 5214 -1648
rect 5180 -1716 5214 -1682
rect 5180 -1750 5214 -1716
rect 5180 -1784 5214 -1750
rect 5180 -1818 5214 -1784
rect 5180 -1852 5214 -1818
rect 5180 -1886 5214 -1852
rect 5180 -1920 5214 -1886
rect 5180 -1954 5214 -1920
rect 5180 -1988 5214 -1954
rect 5180 -2022 5214 -1988
rect 5180 -2056 5214 -2022
rect 5180 -2090 5214 -2056
rect 5180 -2124 5214 -2090
rect 5180 -2158 5214 -2124
rect 5180 -2192 5214 -2158
rect 5180 -2226 5214 -2192
rect 5180 -2260 5214 -2226
rect 5180 -2276 5214 -2260
rect 1934 -2574 1968 -2528
rect 1934 -2608 1968 -2574
rect 1934 -2642 1968 -2608
rect 1934 -2676 1968 -2642
rect 1934 -2710 1968 -2676
rect 1934 -2744 1968 -2710
rect 1934 -2778 1968 -2744
rect 1934 -2812 1968 -2778
rect 1934 -2846 1968 -2812
rect 1934 -2880 1968 -2846
rect 1934 -2914 1968 -2880
rect 1934 -2948 1968 -2914
rect 1934 -2982 1968 -2948
rect 1934 -3016 1968 -2982
rect 1934 -3050 1968 -3016
rect 1934 -3084 1968 -3050
rect 1934 -3118 1968 -3084
rect 1934 -3152 1968 -3118
rect 1934 -3186 1968 -3152
rect 1934 -3220 1968 -3186
rect 1934 -3254 1968 -3220
rect 1934 -3288 1968 -3254
rect 1934 -3304 1968 -3288
rect 3558 -2574 3592 -2528
rect 3558 -2608 3592 -2574
rect 3558 -2642 3592 -2608
rect 3558 -2676 3592 -2642
rect 3558 -2710 3592 -2676
rect 3558 -2744 3592 -2710
rect 3558 -2778 3592 -2744
rect 3558 -2812 3592 -2778
rect 3558 -2846 3592 -2812
rect 3558 -2880 3592 -2846
rect 3558 -2914 3592 -2880
rect 3558 -2948 3592 -2914
rect 3558 -2982 3592 -2948
rect 3558 -3016 3592 -2982
rect 3558 -3050 3592 -3016
rect 3558 -3084 3592 -3050
rect 3558 -3118 3592 -3084
rect 3558 -3152 3592 -3118
rect 3558 -3186 3592 -3152
rect 3558 -3220 3592 -3186
rect 3558 -3254 3592 -3220
rect 3558 -3288 3592 -3254
rect 3558 -3304 3592 -3288
rect 5180 -2574 5214 -2528
rect 5180 -2608 5214 -2574
rect 5180 -2642 5214 -2608
rect 5180 -2676 5214 -2642
rect 5180 -2710 5214 -2676
rect 5180 -2744 5214 -2710
rect 5180 -2778 5214 -2744
rect 5180 -2812 5214 -2778
rect 5180 -2846 5214 -2812
rect 5180 -2880 5214 -2846
rect 5180 -2914 5214 -2880
rect 5180 -2948 5214 -2914
rect 5180 -2982 5214 -2948
rect 5180 -3016 5214 -2982
rect 5180 -3050 5214 -3016
rect 5180 -3084 5214 -3050
rect 5180 -3118 5214 -3084
rect 5180 -3152 5214 -3118
rect 5180 -3186 5214 -3152
rect 5180 -3220 5214 -3186
rect 5180 -3254 5214 -3220
rect 5180 -3288 5214 -3254
rect 5180 -3304 5214 -3288
rect 1933 -3592 1967 -3558
rect 1933 -3626 1967 -3592
rect 1933 -3660 1967 -3626
rect 1933 -3694 1967 -3660
rect 1933 -3728 1967 -3694
rect 1933 -3762 1967 -3728
rect 1933 -3796 1967 -3762
rect 1933 -3830 1967 -3796
rect 1933 -3864 1967 -3830
rect 1933 -3898 1967 -3864
rect 1933 -3932 1967 -3898
rect 1933 -3966 1967 -3932
rect 1933 -4000 1967 -3966
rect 1933 -4034 1967 -4000
rect 1933 -4068 1967 -4034
rect 1933 -4102 1967 -4068
rect 1933 -4136 1967 -4102
rect 1933 -4170 1967 -4136
rect 1933 -4204 1967 -4170
rect 1933 -4238 1967 -4204
rect 1933 -4272 1967 -4238
rect 1933 -4306 1967 -4272
rect 1933 -4340 1967 -4306
rect 1933 -4374 1967 -4340
rect 1933 -4408 1967 -4374
rect 1933 -4442 1967 -4408
rect 1933 -4476 1967 -4442
rect 1933 -4510 1967 -4476
rect 3535 -3592 3569 -3558
rect 3535 -3626 3569 -3592
rect 3535 -3660 3569 -3626
rect 3535 -3694 3569 -3660
rect 3535 -3728 3569 -3694
rect 3535 -3762 3569 -3728
rect 3535 -3796 3569 -3762
rect 3535 -3830 3569 -3796
rect 3535 -3864 3569 -3830
rect 3535 -3898 3569 -3864
rect 3535 -3932 3569 -3898
rect 3535 -3966 3569 -3932
rect 3535 -4000 3569 -3966
rect 3535 -4034 3569 -4000
rect 3535 -4068 3569 -4034
rect 3535 -4102 3569 -4068
rect 3535 -4136 3569 -4102
rect 3535 -4170 3569 -4136
rect 3535 -4204 3569 -4170
rect 3535 -4238 3569 -4204
rect 3535 -4272 3569 -4238
rect 3535 -4306 3569 -4272
rect 3535 -4340 3569 -4306
rect 3535 -4374 3569 -4340
rect 3535 -4408 3569 -4374
rect 3535 -4442 3569 -4408
rect 3535 -4476 3569 -4442
rect 3535 -4510 3569 -4476
rect 5158 -3592 5192 -3558
rect 5158 -3626 5192 -3592
rect 5158 -3660 5192 -3626
rect 5158 -3694 5192 -3660
rect 5158 -3728 5192 -3694
rect 5158 -3762 5192 -3728
rect 5158 -3796 5192 -3762
rect 5158 -3830 5192 -3796
rect 5158 -3864 5192 -3830
rect 5158 -3898 5192 -3864
rect 5158 -3932 5192 -3898
rect 5158 -3966 5192 -3932
rect 5158 -4000 5192 -3966
rect 5158 -4034 5192 -4000
rect 5158 -4068 5192 -4034
rect 5158 -4102 5192 -4068
rect 5158 -4136 5192 -4102
rect 5158 -4170 5192 -4136
rect 5158 -4204 5192 -4170
rect 5158 -4238 5192 -4204
rect 5158 -4272 5192 -4238
rect 5158 -4306 5192 -4272
rect 5158 -4340 5192 -4306
rect 5158 -4374 5192 -4340
rect 5158 -4408 5192 -4374
rect 5158 -4442 5192 -4408
rect 5158 -4476 5192 -4442
rect 5158 -4510 5192 -4476
<< metal1 >>
rect 1914 582 2030 588
rect 1914 112 2030 234
rect 3538 582 3654 588
rect 3538 112 3654 234
rect 5160 582 5276 588
rect 5160 112 5276 234
rect 1914 100 2044 112
rect 1914 -2276 1934 100
rect 1968 -2276 2044 100
rect 1914 -2288 2044 -2276
rect 1712 -2378 1828 -2372
rect 1510 -3976 1684 -3454
rect 1510 -4092 1558 -3976
rect 1674 -4092 1684 -3976
rect 1510 -4254 1684 -4092
rect 1712 -4190 1828 -2436
rect 2058 -2378 2450 -2374
rect 2058 -2436 2196 -2378
rect 2312 -2436 2450 -2378
rect 2058 -2438 2450 -2436
rect 1712 -4254 1828 -4248
rect 1856 -2528 2006 -2516
rect 1856 -3304 1934 -2528
rect 1968 -3304 2006 -2528
rect 1856 -3316 2006 -3304
rect 2478 -3100 2594 112
rect 3538 100 3672 112
rect 2652 -1760 2912 -1644
rect 2652 -3100 2768 -1760
rect 2478 -3122 2768 -3100
rect 2478 -3180 2566 -3122
rect 2682 -3180 2768 -3122
rect 2478 -3204 2768 -3180
rect 2796 -3088 2912 -1760
rect 2940 -1760 3200 -1644
rect 2940 -3088 3056 -1760
rect 2796 -3204 3056 -3088
rect 3084 -3088 3200 -1760
rect 3228 -1666 3510 -1644
rect 3228 -1724 3312 -1666
rect 3428 -1724 3510 -1666
rect 3228 -1748 3510 -1724
rect 3228 -3088 3344 -1748
rect 3394 -2378 3510 -1748
rect 3538 -2276 3558 100
rect 3592 -2276 3672 100
rect 3538 -2288 3672 -2276
rect 3394 -2442 3510 -2436
rect 3682 -2378 4074 -2374
rect 3682 -2436 3820 -2378
rect 3936 -2436 4074 -2378
rect 3682 -2438 4074 -2436
rect 3084 -3204 3344 -3088
rect 3482 -2528 3630 -2516
rect 2478 -3316 2594 -3204
rect 1856 -3546 1972 -3316
rect 2500 -3462 2594 -3316
rect 3482 -3304 3558 -2528
rect 3592 -3304 3630 -2528
rect 3482 -3316 3630 -3304
rect 4102 -3100 4218 112
rect 5160 100 5294 112
rect 4272 -1760 4532 -1644
rect 4272 -3100 4388 -1760
rect 4102 -3122 4388 -3100
rect 4102 -3180 4188 -3122
rect 4304 -3180 4388 -3122
rect 4102 -3204 4388 -3180
rect 4416 -3088 4532 -1760
rect 4560 -1760 4820 -1644
rect 4560 -3088 4676 -1760
rect 4416 -3204 4676 -3088
rect 4704 -3088 4820 -1760
rect 4848 -1666 5132 -1644
rect 4848 -1724 4932 -1666
rect 5048 -1724 5132 -1666
rect 4848 -1748 5132 -1724
rect 4848 -3088 4964 -1748
rect 5016 -2378 5132 -1748
rect 5160 -2276 5180 100
rect 5214 -2276 5294 100
rect 5160 -2288 5294 -2276
rect 5724 -2344 5840 112
rect 6628 -2344 6802 -2054
rect 5016 -2442 5132 -2436
rect 5248 -2375 5306 -2344
rect 5724 -2374 5920 -2344
rect 5248 -2378 5696 -2375
rect 5248 -2436 5442 -2378
rect 5558 -2436 5696 -2378
rect 5248 -2438 5696 -2436
rect 5724 -2432 5804 -2374
rect 5248 -2460 5306 -2438
rect 5724 -2460 5920 -2432
rect 6484 -2374 6802 -2344
rect 6600 -2432 6802 -2374
rect 6484 -2460 6802 -2432
rect 4704 -3204 4964 -3088
rect 5102 -2528 5252 -2516
rect 4102 -3316 4218 -3204
rect 1856 -3558 1973 -3546
rect 1856 -4510 1933 -3558
rect 1967 -4510 1973 -3558
rect 1856 -4522 1973 -4510
rect 1856 -4694 1972 -4522
rect 2517 -4570 2749 -3496
rect 3482 -3558 3598 -3316
rect 4120 -3462 4218 -3316
rect 5102 -3304 5180 -2528
rect 5214 -3304 5252 -2528
rect 5102 -3316 5252 -3304
rect 5724 -3316 5840 -2460
rect 3119 -3974 3189 -3968
rect 3119 -4090 3125 -3974
rect 3183 -4090 3189 -3974
rect 3119 -4096 3189 -4090
rect 3482 -4510 3535 -3558
rect 3569 -4510 3598 -3558
rect 1856 -5048 1972 -5042
rect 3482 -4694 3598 -4510
rect 4120 -4570 4352 -3496
rect 5102 -3546 5218 -3316
rect 5746 -3462 5840 -3316
rect 5102 -3558 5219 -3546
rect 4722 -3974 4792 -3968
rect 4722 -4090 4728 -3974
rect 4786 -4090 4792 -3974
rect 4722 -4096 4792 -4090
rect 5102 -4510 5158 -3558
rect 5192 -4510 5219 -3558
rect 5102 -4522 5219 -4510
rect 3482 -5048 3598 -5042
rect 5102 -4694 5218 -4522
rect 5746 -4570 5978 -3496
rect 6350 -3976 6414 -3970
rect 6408 -4092 6414 -3976
rect 6350 -4098 6414 -4092
rect 6484 -4190 6600 -2460
rect 6628 -2750 6802 -2460
rect 6484 -4254 6600 -4248
rect 5102 -5048 5218 -5042
<< via1 >>
rect 1914 234 2030 582
rect 3538 234 3654 582
rect 5160 234 5276 582
rect 1712 -2436 1828 -2378
rect 1558 -4092 1674 -3976
rect 2196 -2436 2312 -2378
rect 1712 -4248 1828 -4190
rect 2566 -3180 2682 -3122
rect 3312 -1724 3428 -1666
rect 3394 -2436 3510 -2378
rect 3820 -2436 3936 -2378
rect 4188 -3180 4304 -3122
rect 4932 -1724 5048 -1666
rect 5016 -2436 5132 -2378
rect 5442 -2436 5558 -2378
rect 5804 -2432 5920 -2374
rect 6484 -2432 6600 -2374
rect 3125 -4090 3183 -3974
rect 1856 -5042 1972 -4694
rect 4728 -4090 4786 -3974
rect 3482 -5042 3598 -4694
rect 6350 -4092 6408 -3976
rect 6484 -4248 6600 -4190
rect 5102 -5042 5218 -4694
<< metal2 >>
rect 1510 582 6802 690
rect 1510 234 1914 582
rect 2030 234 3538 582
rect 3654 234 5160 582
rect 5276 234 6802 582
rect 1510 222 6802 234
rect 3306 -1666 3434 -1644
rect 3306 -1724 3312 -1666
rect 3428 -1724 3434 -1666
rect 3306 -1748 3434 -1724
rect 4926 -1666 5054 -1644
rect 4926 -1724 4932 -1666
rect 5048 -1724 5054 -1666
rect 4926 -1748 5054 -1724
rect 1712 -2378 2312 -2354
rect 1828 -2436 2196 -2378
rect 1712 -2458 2312 -2436
rect 3394 -2378 3936 -2354
rect 3510 -2436 3820 -2378
rect 3394 -2458 3936 -2436
rect 5016 -2378 5558 -2354
rect 5132 -2436 5442 -2378
rect 5016 -2458 5558 -2436
rect 5782 -2374 6600 -2344
rect 5782 -2432 5804 -2374
rect 5920 -2432 6484 -2374
rect 5782 -2460 6600 -2432
rect 2560 -3122 2688 -3100
rect 2560 -3180 2566 -3122
rect 2682 -3180 2688 -3122
rect 2560 -3204 2688 -3180
rect 4182 -3122 4310 -3100
rect 4182 -3180 4188 -3122
rect 4304 -3180 4310 -3122
rect 4182 -3204 4310 -3180
rect 1552 -3974 6414 -3930
rect 1552 -3976 3125 -3974
rect 1552 -4092 1558 -3976
rect 1674 -4090 3125 -3976
rect 3183 -4090 4728 -3974
rect 4786 -3976 6414 -3974
rect 4786 -4090 6350 -3976
rect 1674 -4092 6350 -4090
rect 6408 -4092 6414 -3976
rect 1552 -4138 6414 -4092
rect 1712 -4190 6600 -4166
rect 1828 -4248 6484 -4190
rect 1712 -4270 6600 -4248
rect 1510 -4694 6802 -4682
rect 1510 -5042 1856 -4694
rect 1972 -5042 3482 -4694
rect 3598 -5042 5102 -4694
rect 5218 -5042 6802 -4694
rect 1510 -5150 6802 -5042
use sky130_fd_pr__pfet_01v8_lvt_5L5ME6  M1
timestamp 1680254034
transform 1 0 2254 0 1 -1088
box -294 -1300 294 1300
use sky130_fd_pr__nfet_01v8_lvt_D8FT7U  M2
timestamp 1680262531
transform 1 0 2254 0 1 -2916
box -258 -488 258 488
use sky130_fd_pr__pfet_01v8_lvt_5L5ME6  M3
timestamp 1680254034
transform 1 0 3878 0 1 -1088
box -294 -1300 294 1300
use sky130_fd_pr__nfet_01v8_lvt_D8FT7U  M4
timestamp 1680262531
transform 1 0 3878 0 1 -2916
box -258 -488 258 488
use sky130_fd_pr__pfet_01v8_lvt_5L5ME6  M5
timestamp 1680254034
transform 1 0 5500 0 1 -1088
box -294 -1300 294 1300
use sky130_fd_pr__nfet_01v8_lvt_D8FT7U  M6
timestamp 1680262531
transform 1 0 5500 0 1 -2916
box -258 -488 258 488
use sky130_fd_pr__cap_var_lvt_SC9F2N  XC1
timestamp 1680254065
transform 1 0 5865 0 1 -4034
box -633 -591 633 591
use sky130_fd_pr__cap_var_lvt_SC9F2N  XC2
timestamp 1680254065
transform 1 0 4244 0 1 -4034
box -633 -591 633 591
use sky130_fd_pr__cap_var_lvt_SC9F2N  XC3
timestamp 1680254065
transform 1 0 2640 0 1 -4034
box -633 -591 633 591
<< labels >>
flabel metal1 6628 -2750 6802 -2054 0 FreeMono 960 90 0 0 vosc
port 3 nsew
flabel metal2 1510 222 6802 690 0 FreeMono 1600 0 0 0 vdd
port 2 nsew
flabel metal2 1510 -5150 6802 -4682 1 FreeMono 1600 0 0 0 vss
port 1 n
flabel metal1 1510 -4254 1684 -3454 0 FreeMono 800 90 0 0 vtemp
port 0 nsew
<< end >>
