magic
tech sky130A
magscale 1 2
timestamp 1681062556
<< error_p >>
rect -29 541 29 547
rect -29 507 -17 541
rect -29 501 29 507
rect -76 -531 -18 469
rect 18 -531 76 469
<< nmoslvt >>
rect -18 -531 18 469
<< ndiff >>
rect -76 457 -18 469
rect -76 -519 -64 457
rect -30 -519 -18 457
rect -76 -531 -18 -519
rect 18 457 76 469
rect 18 -519 30 457
rect 64 -519 76 457
rect 18 -531 76 -519
<< ndiffc >>
rect -64 -519 -30 457
rect 30 -519 64 457
<< poly >>
rect -33 541 33 557
rect -33 507 -17 541
rect 17 507 33 541
rect -33 491 33 507
rect -18 469 18 491
rect -18 -557 18 -531
<< polycont >>
rect -17 507 17 541
<< locali >>
rect -33 507 -17 541
rect 17 507 33 541
rect -64 457 -30 473
rect -64 -535 -30 -519
rect 30 457 64 473
rect 30 -535 64 -519
<< viali >>
rect -17 507 17 541
rect -64 -519 -30 457
rect 30 -519 64 457
<< metal1 >>
rect -29 541 29 547
rect -29 507 -17 541
rect 17 507 29 541
rect -29 501 29 507
rect -70 457 -24 469
rect -70 -519 -64 457
rect -30 -519 -24 457
rect -70 -531 -24 -519
rect 24 457 70 469
rect 24 -519 30 457
rect 64 -519 70 457
rect 24 -531 70 -519
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.0 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
