magic
tech sky130A
magscale 1 2
timestamp 1681321933
<< xpolycontact >>
rect -573 1146 573 1578
rect -573 -1578 573 -1146
<< xpolyres >>
rect -573 -1146 573 1146
<< viali >>
rect -557 1163 557 1560
rect -557 -1560 557 -1163
<< metal1 >>
rect -569 1560 569 1566
rect -569 1163 -557 1560
rect 557 1163 569 1560
rect -569 1157 569 1163
rect -569 -1163 569 -1157
rect -569 -1560 -557 -1163
rect 557 -1560 569 -1163
rect -569 -1566 569 -1560
<< res5p73 >>
rect -575 -1148 575 1148
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 11.46 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 4.065k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
