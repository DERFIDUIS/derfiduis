magic
tech sky130A
magscale 1 2
timestamp 1680265380
<< metal3 >>
rect -3186 6172 3186 6200
rect -3186 148 3102 6172
rect 3166 148 3186 6172
rect -3186 120 3186 148
rect -3186 -148 3186 -120
rect -3186 -6172 3102 -148
rect 3166 -6172 3186 -148
rect -3186 -6200 3186 -6172
<< via3 >>
rect 3102 148 3166 6172
rect 3102 -6172 3166 -148
<< mimcap >>
rect -3146 6120 2854 6160
rect -3146 200 -3106 6120
rect 2814 200 2854 6120
rect -3146 160 2854 200
rect -3146 -200 2854 -160
rect -3146 -6120 -3106 -200
rect 2814 -6120 2854 -200
rect -3146 -6160 2854 -6120
<< mimcapcontact >>
rect -3106 200 2814 6120
rect -3106 -6120 2814 -200
<< metal4 >>
rect -198 6121 -94 6320
rect 3082 6172 3186 6320
rect -3107 6120 2815 6121
rect -3107 200 -3106 6120
rect 2814 200 2815 6120
rect -3107 199 2815 200
rect -198 -199 -94 199
rect 3082 148 3102 6172
rect 3166 148 3186 6172
rect 3082 -148 3186 148
rect -3107 -200 2815 -199
rect -3107 -6120 -3106 -200
rect 2814 -6120 2815 -200
rect -3107 -6121 2815 -6120
rect -198 -6320 -94 -6121
rect 3082 -6172 3102 -148
rect 3166 -6172 3186 -148
rect 3082 -6320 3186 -6172
<< properties >>
string FIXED_BBOX -3186 120 2894 6200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 30.0 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
