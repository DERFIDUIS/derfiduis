magic
tech sky130A
magscale 1 2
timestamp 1682114810
<< nwell >>
rect -5328 -1526 -5170 -1432
rect -5328 -1528 -5164 -1526
rect -5334 -1994 -5164 -1528
rect -4396 -1994 -4254 -1432
rect -5334 -2258 -5198 -2248
rect -5300 -2310 -5164 -2258
rect -5298 -2348 -5164 -2310
rect -5334 -2810 -5164 -2348
rect -340 -2302 -224 -1246
rect -340 -2408 -174 -2302
rect 726 -2408 840 -1246
rect 1790 -2408 1904 -1246
rect 2854 -2408 2968 -1246
rect 3930 -2408 4034 -1246
<< nbase >>
rect -2770 -4238 -2742 -4198
rect -2480 -4204 -2466 -4198
rect -2486 -4238 -2466 -4204
rect -1630 -4214 -1622 -4178
rect -1574 -4238 -1556 -4204
rect -2766 -4274 -2762 -4238
rect -2770 -4406 -2726 -4274
rect -2766 -4414 -2762 -4406
rect -2766 -4482 -2760 -4414
rect -2480 -4482 -2472 -4238
rect -1572 -4274 -1568 -4238
rect -1578 -4406 -1558 -4274
rect -1572 -4474 -1568 -4406
rect -1572 -4482 -1566 -4474
rect -1290 -4482 -1284 -4474
rect -2766 -4488 -2474 -4482
rect -1572 -4488 -1284 -4482
<< ndiff >>
rect -3158 -2108 -3156 -1308
rect -3070 -2108 -3068 -1308
rect -2094 -2108 -2092 -1308
rect -2006 -2108 -2004 -1308
rect -1030 -2108 -1028 -1308
rect -942 -2108 -940 -1308
rect -5294 -3060 -5292 -2960
rect -5206 -3060 -5204 -2960
rect -3070 -3662 -3068 -2862
rect -2094 -3662 -2092 -2862
rect -2006 -3662 -2004 -2862
rect -1030 -3662 -1028 -2862
rect -942 -3662 -940 -2862
rect 62 -3136 64 -2936
rect 438 -3136 440 -2936
rect 526 -3136 528 -2936
rect 1502 -3136 1504 -2936
rect 2190 -3136 2192 -2936
rect 2566 -3136 2568 -2936
rect 2654 -3136 2656 -2936
rect 3630 -3136 3632 -2936
rect 1264 -4880 1266 -3880
rect 1352 -4880 1354 -3880
rect 2328 -4880 2330 -3880
rect 2416 -4880 2418 -3880
<< pdiff >>
rect -5294 -1932 -5292 -1532
rect -5206 -1932 -5204 -1532
rect -4296 -1894 -4294 -1494
rect -238 -2308 -236 -1308
rect 738 -2308 740 -1308
rect 826 -2308 828 -1308
rect 1802 -2308 1804 -1308
rect 1890 -2308 1892 -1308
rect 2866 -2308 2868 -1308
rect 2954 -2308 2956 -1308
rect 3930 -2308 3932 -1308
rect -5294 -2748 -5292 -2348
rect -5206 -2748 -5204 -2348
<< psubdiff >>
rect -3156 -1366 -3070 -1308
rect -3156 -1400 -3130 -1366
rect -3096 -1400 -3070 -1366
rect -3156 -1434 -3070 -1400
rect -3156 -1468 -3130 -1434
rect -3096 -1468 -3070 -1434
rect -3156 -1502 -3070 -1468
rect -3156 -1536 -3130 -1502
rect -3096 -1536 -3070 -1502
rect -3156 -1570 -3070 -1536
rect -3156 -1604 -3130 -1570
rect -3096 -1604 -3070 -1570
rect -3156 -1638 -3070 -1604
rect -3156 -1672 -3130 -1638
rect -3096 -1672 -3070 -1638
rect -3156 -1706 -3070 -1672
rect -3156 -1740 -3130 -1706
rect -3096 -1740 -3070 -1706
rect -3156 -1774 -3070 -1740
rect -3156 -1808 -3130 -1774
rect -3096 -1808 -3070 -1774
rect -3156 -1842 -3070 -1808
rect -3156 -1876 -3130 -1842
rect -3096 -1876 -3070 -1842
rect -3156 -1910 -3070 -1876
rect -3156 -1944 -3130 -1910
rect -3096 -1944 -3070 -1910
rect -3156 -1978 -3070 -1944
rect -3156 -2012 -3130 -1978
rect -3096 -2012 -3070 -1978
rect -3156 -2046 -3070 -2012
rect -3156 -2080 -3130 -2046
rect -3096 -2080 -3070 -2046
rect -3156 -2108 -3070 -2080
rect -2092 -1366 -2006 -1308
rect -2092 -1400 -2066 -1366
rect -2032 -1400 -2006 -1366
rect -2092 -1434 -2006 -1400
rect -2092 -1468 -2066 -1434
rect -2032 -1468 -2006 -1434
rect -2092 -1502 -2006 -1468
rect -2092 -1536 -2066 -1502
rect -2032 -1536 -2006 -1502
rect -2092 -1570 -2006 -1536
rect -2092 -1604 -2066 -1570
rect -2032 -1604 -2006 -1570
rect -2092 -1638 -2006 -1604
rect -2092 -1672 -2066 -1638
rect -2032 -1672 -2006 -1638
rect -2092 -1706 -2006 -1672
rect -2092 -1740 -2066 -1706
rect -2032 -1740 -2006 -1706
rect -2092 -1774 -2006 -1740
rect -2092 -1808 -2066 -1774
rect -2032 -1808 -2006 -1774
rect -2092 -1842 -2006 -1808
rect -2092 -1876 -2066 -1842
rect -2032 -1876 -2006 -1842
rect -2092 -1910 -2006 -1876
rect -2092 -1944 -2066 -1910
rect -2032 -1944 -2006 -1910
rect -2092 -1978 -2006 -1944
rect -2092 -2012 -2066 -1978
rect -2032 -2012 -2006 -1978
rect -2092 -2046 -2006 -2012
rect -2092 -2080 -2066 -2046
rect -2032 -2080 -2006 -2046
rect -2092 -2108 -2006 -2080
rect -1028 -1366 -942 -1308
rect -1028 -1400 -1002 -1366
rect -968 -1400 -942 -1366
rect -1028 -1434 -942 -1400
rect -1028 -1468 -1002 -1434
rect -968 -1468 -942 -1434
rect -1028 -1502 -942 -1468
rect -1028 -1536 -1002 -1502
rect -968 -1536 -942 -1502
rect -1028 -1570 -942 -1536
rect -1028 -1604 -1002 -1570
rect -968 -1604 -942 -1570
rect -1028 -1638 -942 -1604
rect -1028 -1672 -1002 -1638
rect -968 -1672 -942 -1638
rect -1028 -1706 -942 -1672
rect -1028 -1740 -1002 -1706
rect -968 -1740 -942 -1706
rect -1028 -1774 -942 -1740
rect -1028 -1808 -1002 -1774
rect -968 -1808 -942 -1774
rect -1028 -1842 -942 -1808
rect -1028 -1876 -1002 -1842
rect -968 -1876 -942 -1842
rect -1028 -1910 -942 -1876
rect -1028 -1944 -1002 -1910
rect -968 -1944 -942 -1910
rect -1028 -1978 -942 -1944
rect -1028 -2012 -1002 -1978
rect -968 -2012 -942 -1978
rect -1028 -2046 -942 -2012
rect -1028 -2080 -1002 -2046
rect -968 -2080 -942 -2046
rect -1028 -2108 -942 -2080
rect -3134 -2920 -3070 -2862
rect -3134 -2954 -3130 -2920
rect -3096 -2954 -3070 -2920
rect -5292 -2986 -5206 -2960
rect -5292 -3032 -5266 -2986
rect -5232 -3032 -5206 -2986
rect -5292 -3060 -5206 -3032
rect -3134 -2988 -3070 -2954
rect -3134 -3022 -3130 -2988
rect -3096 -3022 -3070 -2988
rect -3134 -3056 -3070 -3022
rect -3134 -3090 -3130 -3056
rect -3096 -3090 -3070 -3056
rect -3134 -3124 -3070 -3090
rect -3134 -3158 -3130 -3124
rect -3096 -3158 -3070 -3124
rect -3134 -3192 -3070 -3158
rect -3134 -3226 -3130 -3192
rect -3096 -3226 -3070 -3192
rect -3134 -3260 -3070 -3226
rect -3134 -3294 -3130 -3260
rect -3096 -3294 -3070 -3260
rect -3134 -3328 -3070 -3294
rect -3134 -3362 -3130 -3328
rect -3096 -3362 -3070 -3328
rect -3134 -3396 -3070 -3362
rect -3134 -3430 -3130 -3396
rect -3096 -3430 -3070 -3396
rect -3134 -3464 -3070 -3430
rect -3134 -3498 -3130 -3464
rect -3096 -3498 -3070 -3464
rect -3134 -3532 -3070 -3498
rect -3134 -3566 -3130 -3532
rect -3096 -3566 -3070 -3532
rect -3134 -3600 -3070 -3566
rect -3134 -3634 -3130 -3600
rect -3096 -3634 -3070 -3600
rect -3134 -3662 -3070 -3634
rect -2092 -2920 -2006 -2862
rect -2092 -2954 -2066 -2920
rect -2032 -2954 -2006 -2920
rect -2092 -2988 -2006 -2954
rect -2092 -3022 -2066 -2988
rect -2032 -3022 -2006 -2988
rect -2092 -3056 -2006 -3022
rect -2092 -3090 -2066 -3056
rect -2032 -3090 -2006 -3056
rect -2092 -3124 -2006 -3090
rect -2092 -3158 -2066 -3124
rect -2032 -3158 -2006 -3124
rect -2092 -3192 -2006 -3158
rect -2092 -3226 -2066 -3192
rect -2032 -3226 -2006 -3192
rect -2092 -3260 -2006 -3226
rect -2092 -3294 -2066 -3260
rect -2032 -3294 -2006 -3260
rect -2092 -3328 -2006 -3294
rect -2092 -3362 -2066 -3328
rect -2032 -3362 -2006 -3328
rect -2092 -3396 -2006 -3362
rect -2092 -3430 -2066 -3396
rect -2032 -3430 -2006 -3396
rect -2092 -3464 -2006 -3430
rect -2092 -3498 -2066 -3464
rect -2032 -3498 -2006 -3464
rect -2092 -3532 -2006 -3498
rect -2092 -3566 -2066 -3532
rect -2032 -3566 -2006 -3532
rect -2092 -3600 -2006 -3566
rect -2092 -3634 -2066 -3600
rect -2032 -3634 -2006 -3600
rect -2092 -3662 -2006 -3634
rect -1028 -2920 -942 -2862
rect -1028 -2954 -1002 -2920
rect -968 -2954 -942 -2920
rect -1028 -2988 -942 -2954
rect -1028 -3022 -1002 -2988
rect -968 -3022 -942 -2988
rect -1028 -3056 -942 -3022
rect -1028 -3090 -1002 -3056
rect -968 -3090 -942 -3056
rect -1028 -3124 -942 -3090
rect -1028 -3158 -1002 -3124
rect -968 -3158 -942 -3124
rect -1028 -3192 -942 -3158
rect -1028 -3226 -1002 -3192
rect -968 -3226 -942 -3192
rect -1028 -3260 -942 -3226
rect -1028 -3294 -1002 -3260
rect -968 -3294 -942 -3260
rect -1028 -3328 -942 -3294
rect -1028 -3362 -1002 -3328
rect -968 -3362 -942 -3328
rect -1028 -3396 -942 -3362
rect -1028 -3430 -1002 -3396
rect -968 -3430 -942 -3396
rect -1028 -3464 -942 -3430
rect -1028 -3498 -1002 -3464
rect -968 -3498 -942 -3464
rect -1028 -3532 -942 -3498
rect -1028 -3566 -1002 -3532
rect -968 -3566 -942 -3532
rect -1028 -3600 -942 -3566
rect -1028 -3634 -1002 -3600
rect -968 -3634 -942 -3600
rect -1028 -3662 -942 -3634
rect -2 -2990 62 -2936
rect -2 -3024 2 -2990
rect 36 -3024 62 -2990
rect -2 -3058 62 -3024
rect -2 -3092 2 -3058
rect 36 -3092 62 -3058
rect -2 -3136 62 -3092
rect 440 -2990 526 -2936
rect 440 -3024 466 -2990
rect 500 -3024 526 -2990
rect 440 -3058 526 -3024
rect 440 -3092 466 -3058
rect 500 -3092 526 -3058
rect 440 -3136 526 -3092
rect 1504 -2990 1568 -2936
rect 1504 -3024 1530 -2990
rect 1564 -3024 1568 -2990
rect 1504 -3058 1568 -3024
rect 1504 -3092 1530 -3058
rect 1564 -3092 1568 -3058
rect 1504 -3136 1568 -3092
rect 2126 -2990 2190 -2936
rect 2126 -3024 2130 -2990
rect 2164 -3024 2190 -2990
rect 2126 -3058 2190 -3024
rect 2126 -3092 2130 -3058
rect 2164 -3092 2190 -3058
rect 2126 -3136 2190 -3092
rect 2568 -2990 2654 -2936
rect 2568 -3024 2594 -2990
rect 2628 -3024 2654 -2990
rect 2568 -3058 2654 -3024
rect 2568 -3092 2594 -3058
rect 2628 -3092 2654 -3058
rect 2568 -3136 2654 -3092
rect 3632 -2990 3696 -2936
rect 3632 -3024 3658 -2990
rect 3692 -3024 3696 -2990
rect 3632 -3058 3696 -3024
rect 3632 -3092 3658 -3058
rect 3692 -3092 3696 -3058
rect 3632 -3136 3696 -3092
rect 1266 -3934 1352 -3880
rect 1266 -3968 1292 -3934
rect 1326 -3968 1352 -3934
rect 1266 -4002 1352 -3968
rect 1266 -4036 1292 -4002
rect 1326 -4036 1352 -4002
rect 1266 -4070 1352 -4036
rect 1266 -4104 1292 -4070
rect 1326 -4104 1352 -4070
rect 1266 -4138 1352 -4104
rect 1266 -4172 1292 -4138
rect 1326 -4172 1352 -4138
rect 1266 -4206 1352 -4172
rect 1266 -4240 1292 -4206
rect 1326 -4240 1352 -4206
rect 1266 -4274 1352 -4240
rect 1266 -4308 1292 -4274
rect 1326 -4308 1352 -4274
rect 1266 -4342 1352 -4308
rect 1266 -4376 1292 -4342
rect 1326 -4376 1352 -4342
rect 1266 -4410 1352 -4376
rect 1266 -4444 1292 -4410
rect 1326 -4444 1352 -4410
rect 1266 -4478 1352 -4444
rect 1266 -4512 1292 -4478
rect 1326 -4512 1352 -4478
rect 1266 -4546 1352 -4512
rect 1266 -4580 1292 -4546
rect 1326 -4580 1352 -4546
rect 1266 -4614 1352 -4580
rect 1266 -4648 1292 -4614
rect 1326 -4648 1352 -4614
rect 1266 -4682 1352 -4648
rect 1266 -4716 1292 -4682
rect 1326 -4716 1352 -4682
rect 1266 -4750 1352 -4716
rect 1266 -4784 1292 -4750
rect 1326 -4784 1352 -4750
rect 1266 -4818 1352 -4784
rect 1266 -4852 1292 -4818
rect 1326 -4852 1352 -4818
rect 1266 -4880 1352 -4852
rect 2330 -3934 2416 -3880
rect 2330 -3968 2356 -3934
rect 2390 -3968 2416 -3934
rect 2330 -4002 2416 -3968
rect 2330 -4036 2356 -4002
rect 2390 -4036 2416 -4002
rect 2330 -4070 2416 -4036
rect 2330 -4104 2356 -4070
rect 2390 -4104 2416 -4070
rect 2330 -4138 2416 -4104
rect 2330 -4172 2356 -4138
rect 2390 -4172 2416 -4138
rect 2330 -4206 2416 -4172
rect 2330 -4240 2356 -4206
rect 2390 -4240 2416 -4206
rect 2330 -4274 2416 -4240
rect 2330 -4308 2356 -4274
rect 2390 -4308 2416 -4274
rect 2330 -4342 2416 -4308
rect 2330 -4376 2356 -4342
rect 2390 -4376 2416 -4342
rect 2330 -4410 2416 -4376
rect 2330 -4444 2356 -4410
rect 2390 -4444 2416 -4410
rect 2330 -4478 2416 -4444
rect 2330 -4512 2356 -4478
rect 2390 -4512 2416 -4478
rect 2330 -4546 2416 -4512
rect 2330 -4580 2356 -4546
rect 2390 -4580 2416 -4546
rect 2330 -4614 2416 -4580
rect 2330 -4648 2356 -4614
rect 2390 -4648 2416 -4614
rect 2330 -4682 2416 -4648
rect 2330 -4716 2356 -4682
rect 2390 -4716 2416 -4682
rect 2330 -4750 2416 -4716
rect 2330 -4784 2356 -4750
rect 2390 -4784 2416 -4750
rect 2330 -4818 2416 -4784
rect 2330 -4852 2356 -4818
rect 2390 -4852 2416 -4818
rect 2330 -4880 2416 -4852
<< nsubdiff >>
rect -5292 -1560 -5206 -1532
rect -5292 -1594 -5266 -1560
rect -5232 -1594 -5206 -1560
rect -5292 -1628 -5206 -1594
rect -5292 -1662 -5266 -1628
rect -5232 -1662 -5206 -1628
rect -5292 -1696 -5206 -1662
rect -5292 -1730 -5266 -1696
rect -5232 -1730 -5206 -1696
rect -5292 -1764 -5206 -1730
rect -5292 -1798 -5266 -1764
rect -5232 -1798 -5206 -1764
rect -5292 -1832 -5206 -1798
rect -5292 -1866 -5266 -1832
rect -5232 -1866 -5206 -1832
rect -5292 -1932 -5206 -1866
rect -4360 -1560 -4296 -1494
rect -4360 -1594 -4356 -1560
rect -4322 -1594 -4296 -1560
rect -4360 -1628 -4296 -1594
rect -4360 -1662 -4356 -1628
rect -4322 -1662 -4296 -1628
rect -4360 -1696 -4296 -1662
rect -4360 -1730 -4356 -1696
rect -4322 -1730 -4296 -1696
rect -4360 -1764 -4296 -1730
rect -4360 -1798 -4356 -1764
rect -4322 -1798 -4296 -1764
rect -4360 -1832 -4296 -1798
rect -4360 -1866 -4356 -1832
rect -4322 -1866 -4296 -1832
rect -4360 -1894 -4296 -1866
rect -304 -1362 -238 -1308
rect -304 -1396 -298 -1362
rect -264 -1396 -238 -1362
rect -304 -1430 -238 -1396
rect -304 -1464 -298 -1430
rect -264 -1464 -238 -1430
rect -304 -1498 -238 -1464
rect -304 -1532 -298 -1498
rect -264 -1532 -238 -1498
rect -304 -1566 -238 -1532
rect -304 -1600 -298 -1566
rect -264 -1600 -238 -1566
rect -304 -1634 -238 -1600
rect -304 -1668 -298 -1634
rect -264 -1668 -238 -1634
rect -304 -1702 -238 -1668
rect -304 -1736 -298 -1702
rect -264 -1736 -238 -1702
rect -304 -1770 -238 -1736
rect -304 -1804 -298 -1770
rect -264 -1804 -238 -1770
rect -304 -1838 -238 -1804
rect -304 -1872 -298 -1838
rect -264 -1872 -238 -1838
rect -304 -1906 -238 -1872
rect -304 -1940 -298 -1906
rect -264 -1940 -238 -1906
rect -304 -1974 -238 -1940
rect -304 -2008 -298 -1974
rect -264 -2008 -238 -1974
rect -304 -2042 -238 -2008
rect -304 -2076 -298 -2042
rect -264 -2076 -238 -2042
rect -304 -2110 -238 -2076
rect -304 -2144 -298 -2110
rect -264 -2144 -238 -2110
rect -304 -2178 -238 -2144
rect -304 -2212 -298 -2178
rect -264 -2212 -238 -2178
rect -304 -2246 -238 -2212
rect -304 -2280 -298 -2246
rect -264 -2280 -238 -2246
rect -304 -2308 -238 -2280
rect 740 -1362 826 -1308
rect 740 -1396 766 -1362
rect 800 -1396 826 -1362
rect 740 -1430 826 -1396
rect 740 -1464 766 -1430
rect 800 -1464 826 -1430
rect 740 -1498 826 -1464
rect 740 -1532 766 -1498
rect 800 -1532 826 -1498
rect 740 -1566 826 -1532
rect 740 -1600 766 -1566
rect 800 -1600 826 -1566
rect 740 -1634 826 -1600
rect 740 -1668 766 -1634
rect 800 -1668 826 -1634
rect 740 -1702 826 -1668
rect 740 -1736 766 -1702
rect 800 -1736 826 -1702
rect 740 -1770 826 -1736
rect 740 -1804 766 -1770
rect 800 -1804 826 -1770
rect 740 -1838 826 -1804
rect 740 -1872 766 -1838
rect 800 -1872 826 -1838
rect 740 -1906 826 -1872
rect 740 -1940 766 -1906
rect 800 -1940 826 -1906
rect 740 -1974 826 -1940
rect 740 -2008 766 -1974
rect 800 -2008 826 -1974
rect 740 -2042 826 -2008
rect 740 -2076 766 -2042
rect 800 -2076 826 -2042
rect 740 -2110 826 -2076
rect 740 -2144 766 -2110
rect 800 -2144 826 -2110
rect 740 -2178 826 -2144
rect 740 -2212 766 -2178
rect 800 -2212 826 -2178
rect 740 -2246 826 -2212
rect 740 -2280 766 -2246
rect 800 -2280 826 -2246
rect 740 -2308 826 -2280
rect 1804 -1362 1890 -1308
rect 1804 -1396 1830 -1362
rect 1864 -1396 1890 -1362
rect 1804 -1430 1890 -1396
rect 1804 -1464 1830 -1430
rect 1864 -1464 1890 -1430
rect 1804 -1498 1890 -1464
rect 1804 -1532 1830 -1498
rect 1864 -1532 1890 -1498
rect 1804 -1566 1890 -1532
rect 1804 -1600 1830 -1566
rect 1864 -1600 1890 -1566
rect 1804 -1634 1890 -1600
rect 1804 -1668 1830 -1634
rect 1864 -1668 1890 -1634
rect 1804 -1702 1890 -1668
rect 1804 -1736 1830 -1702
rect 1864 -1736 1890 -1702
rect 1804 -1770 1890 -1736
rect 1804 -1804 1830 -1770
rect 1864 -1804 1890 -1770
rect 1804 -1838 1890 -1804
rect 1804 -1872 1830 -1838
rect 1864 -1872 1890 -1838
rect 1804 -1906 1890 -1872
rect 1804 -1940 1830 -1906
rect 1864 -1940 1890 -1906
rect 1804 -1974 1890 -1940
rect 1804 -2008 1830 -1974
rect 1864 -2008 1890 -1974
rect 1804 -2042 1890 -2008
rect 1804 -2076 1830 -2042
rect 1864 -2076 1890 -2042
rect 1804 -2110 1890 -2076
rect 1804 -2144 1830 -2110
rect 1864 -2144 1890 -2110
rect 1804 -2178 1890 -2144
rect 1804 -2212 1830 -2178
rect 1864 -2212 1890 -2178
rect 1804 -2246 1890 -2212
rect 1804 -2280 1830 -2246
rect 1864 -2280 1890 -2246
rect 1804 -2308 1890 -2280
rect 2868 -1362 2954 -1308
rect 2868 -1396 2894 -1362
rect 2928 -1396 2954 -1362
rect 2868 -1430 2954 -1396
rect 2868 -1464 2894 -1430
rect 2928 -1464 2954 -1430
rect 2868 -1498 2954 -1464
rect 2868 -1532 2894 -1498
rect 2928 -1532 2954 -1498
rect 2868 -1566 2954 -1532
rect 2868 -1600 2894 -1566
rect 2928 -1600 2954 -1566
rect 2868 -1634 2954 -1600
rect 2868 -1668 2894 -1634
rect 2928 -1668 2954 -1634
rect 2868 -1702 2954 -1668
rect 2868 -1736 2894 -1702
rect 2928 -1736 2954 -1702
rect 2868 -1770 2954 -1736
rect 2868 -1804 2894 -1770
rect 2928 -1804 2954 -1770
rect 2868 -1838 2954 -1804
rect 2868 -1872 2894 -1838
rect 2928 -1872 2954 -1838
rect 2868 -1906 2954 -1872
rect 2868 -1940 2894 -1906
rect 2928 -1940 2954 -1906
rect 2868 -1974 2954 -1940
rect 2868 -2008 2894 -1974
rect 2928 -2008 2954 -1974
rect 2868 -2042 2954 -2008
rect 2868 -2076 2894 -2042
rect 2928 -2076 2954 -2042
rect 2868 -2110 2954 -2076
rect 2868 -2144 2894 -2110
rect 2928 -2144 2954 -2110
rect 2868 -2178 2954 -2144
rect 2868 -2212 2894 -2178
rect 2928 -2212 2954 -2178
rect 2868 -2246 2954 -2212
rect 2868 -2280 2894 -2246
rect 2928 -2280 2954 -2246
rect 2868 -2308 2954 -2280
rect 3932 -1362 3998 -1308
rect 3932 -1396 3958 -1362
rect 3992 -1396 3998 -1362
rect 3932 -1430 3998 -1396
rect 3932 -1464 3958 -1430
rect 3992 -1464 3998 -1430
rect 3932 -1498 3998 -1464
rect 3932 -1532 3958 -1498
rect 3992 -1532 3998 -1498
rect 3932 -1566 3998 -1532
rect 3932 -1600 3958 -1566
rect 3992 -1600 3998 -1566
rect 3932 -1634 3998 -1600
rect 3932 -1668 3958 -1634
rect 3992 -1668 3998 -1634
rect 3932 -1702 3998 -1668
rect 3932 -1736 3958 -1702
rect 3992 -1736 3998 -1702
rect 3932 -1770 3998 -1736
rect 3932 -1804 3958 -1770
rect 3992 -1804 3998 -1770
rect 3932 -1838 3998 -1804
rect 3932 -1872 3958 -1838
rect 3992 -1872 3998 -1838
rect 3932 -1906 3998 -1872
rect 3932 -1940 3958 -1906
rect 3992 -1940 3998 -1906
rect 3932 -1974 3998 -1940
rect 3932 -2008 3958 -1974
rect 3992 -2008 3998 -1974
rect 3932 -2042 3998 -2008
rect 3932 -2076 3958 -2042
rect 3992 -2076 3998 -2042
rect 3932 -2110 3998 -2076
rect 3932 -2144 3958 -2110
rect 3992 -2144 3998 -2110
rect 3932 -2178 3998 -2144
rect 3932 -2212 3958 -2178
rect 3992 -2212 3998 -2178
rect 3932 -2246 3998 -2212
rect 3932 -2280 3958 -2246
rect 3992 -2280 3998 -2246
rect 3932 -2308 3998 -2280
rect -5292 -2376 -5206 -2348
rect -5292 -2410 -5266 -2376
rect -5232 -2410 -5206 -2376
rect -5292 -2444 -5206 -2410
rect -5292 -2478 -5266 -2444
rect -5232 -2478 -5206 -2444
rect -5292 -2512 -5206 -2478
rect -5292 -2546 -5266 -2512
rect -5232 -2546 -5206 -2512
rect -5292 -2580 -5206 -2546
rect -5292 -2614 -5266 -2580
rect -5232 -2614 -5206 -2580
rect -5292 -2648 -5206 -2614
rect -5292 -2682 -5266 -2648
rect -5232 -2682 -5206 -2648
rect -5292 -2748 -5206 -2682
rect -2766 -4414 -2762 -4198
rect -2766 -4482 -2760 -4414
rect -2480 -4482 -2472 -4198
rect -1630 -4214 -1622 -4178
rect -1572 -4482 -1566 -4474
rect -1290 -4482 -1284 -4474
rect -2766 -4488 -2474 -4482
rect -1572 -4488 -1284 -4482
<< psubdiffcont >>
rect -3130 -1400 -3096 -1366
rect -3130 -1468 -3096 -1434
rect -3130 -1536 -3096 -1502
rect -3130 -1604 -3096 -1570
rect -3130 -1672 -3096 -1638
rect -3130 -1740 -3096 -1706
rect -3130 -1808 -3096 -1774
rect -3130 -1876 -3096 -1842
rect -3130 -1944 -3096 -1910
rect -3130 -2012 -3096 -1978
rect -3130 -2080 -3096 -2046
rect -2066 -1400 -2032 -1366
rect -2066 -1468 -2032 -1434
rect -2066 -1536 -2032 -1502
rect -2066 -1604 -2032 -1570
rect -2066 -1672 -2032 -1638
rect -2066 -1740 -2032 -1706
rect -2066 -1808 -2032 -1774
rect -2066 -1876 -2032 -1842
rect -2066 -1944 -2032 -1910
rect -2066 -2012 -2032 -1978
rect -2066 -2080 -2032 -2046
rect -1002 -1400 -968 -1366
rect -1002 -1468 -968 -1434
rect -1002 -1536 -968 -1502
rect -1002 -1604 -968 -1570
rect -1002 -1672 -968 -1638
rect -1002 -1740 -968 -1706
rect -1002 -1808 -968 -1774
rect -1002 -1876 -968 -1842
rect -1002 -1944 -968 -1910
rect -1002 -2012 -968 -1978
rect -1002 -2080 -968 -2046
rect -3130 -2954 -3096 -2920
rect -5266 -3032 -5232 -2986
rect -3130 -3022 -3096 -2988
rect -3130 -3090 -3096 -3056
rect -3130 -3158 -3096 -3124
rect -3130 -3226 -3096 -3192
rect -3130 -3294 -3096 -3260
rect -3130 -3362 -3096 -3328
rect -3130 -3430 -3096 -3396
rect -3130 -3498 -3096 -3464
rect -3130 -3566 -3096 -3532
rect -3130 -3634 -3096 -3600
rect -2066 -2954 -2032 -2920
rect -2066 -3022 -2032 -2988
rect -2066 -3090 -2032 -3056
rect -2066 -3158 -2032 -3124
rect -2066 -3226 -2032 -3192
rect -2066 -3294 -2032 -3260
rect -2066 -3362 -2032 -3328
rect -2066 -3430 -2032 -3396
rect -2066 -3498 -2032 -3464
rect -2066 -3566 -2032 -3532
rect -2066 -3634 -2032 -3600
rect -1002 -2954 -968 -2920
rect -1002 -3022 -968 -2988
rect -1002 -3090 -968 -3056
rect -1002 -3158 -968 -3124
rect -1002 -3226 -968 -3192
rect -1002 -3294 -968 -3260
rect -1002 -3362 -968 -3328
rect -1002 -3430 -968 -3396
rect -1002 -3498 -968 -3464
rect -1002 -3566 -968 -3532
rect -1002 -3634 -968 -3600
rect 2 -3024 36 -2990
rect 2 -3092 36 -3058
rect 466 -3024 500 -2990
rect 466 -3092 500 -3058
rect 1530 -3024 1564 -2990
rect 1530 -3092 1564 -3058
rect 2130 -3024 2164 -2990
rect 2130 -3092 2164 -3058
rect 2594 -3024 2628 -2990
rect 2594 -3092 2628 -3058
rect 3658 -3024 3692 -2990
rect 3658 -3092 3692 -3058
rect 1292 -3968 1326 -3934
rect 1292 -4036 1326 -4002
rect 1292 -4104 1326 -4070
rect 1292 -4172 1326 -4138
rect 1292 -4240 1326 -4206
rect 1292 -4308 1326 -4274
rect 1292 -4376 1326 -4342
rect 1292 -4444 1326 -4410
rect 1292 -4512 1326 -4478
rect 1292 -4580 1326 -4546
rect 1292 -4648 1326 -4614
rect 1292 -4716 1326 -4682
rect 1292 -4784 1326 -4750
rect 1292 -4852 1326 -4818
rect 2356 -3968 2390 -3934
rect 2356 -4036 2390 -4002
rect 2356 -4104 2390 -4070
rect 2356 -4172 2390 -4138
rect 2356 -4240 2390 -4206
rect 2356 -4308 2390 -4274
rect 2356 -4376 2390 -4342
rect 2356 -4444 2390 -4410
rect 2356 -4512 2390 -4478
rect 2356 -4580 2390 -4546
rect 2356 -4648 2390 -4614
rect 2356 -4716 2390 -4682
rect 2356 -4784 2390 -4750
rect 2356 -4852 2390 -4818
<< nsubdiffcont >>
rect -5266 -1594 -5232 -1560
rect -5266 -1662 -5232 -1628
rect -5266 -1730 -5232 -1696
rect -5266 -1798 -5232 -1764
rect -5266 -1866 -5232 -1832
rect -4356 -1594 -4322 -1560
rect -4356 -1662 -4322 -1628
rect -4356 -1730 -4322 -1696
rect -4356 -1798 -4322 -1764
rect -4356 -1866 -4322 -1832
rect -298 -1396 -264 -1362
rect -298 -1464 -264 -1430
rect -298 -1532 -264 -1498
rect -298 -1600 -264 -1566
rect -298 -1668 -264 -1634
rect -298 -1736 -264 -1702
rect -298 -1804 -264 -1770
rect -298 -1872 -264 -1838
rect -298 -1940 -264 -1906
rect -298 -2008 -264 -1974
rect -298 -2076 -264 -2042
rect -298 -2144 -264 -2110
rect -298 -2212 -264 -2178
rect -298 -2280 -264 -2246
rect 766 -1396 800 -1362
rect 766 -1464 800 -1430
rect 766 -1532 800 -1498
rect 766 -1600 800 -1566
rect 766 -1668 800 -1634
rect 766 -1736 800 -1702
rect 766 -1804 800 -1770
rect 766 -1872 800 -1838
rect 766 -1940 800 -1906
rect 766 -2008 800 -1974
rect 766 -2076 800 -2042
rect 766 -2144 800 -2110
rect 766 -2212 800 -2178
rect 766 -2280 800 -2246
rect 1830 -1396 1864 -1362
rect 1830 -1464 1864 -1430
rect 1830 -1532 1864 -1498
rect 1830 -1600 1864 -1566
rect 1830 -1668 1864 -1634
rect 1830 -1736 1864 -1702
rect 1830 -1804 1864 -1770
rect 1830 -1872 1864 -1838
rect 1830 -1940 1864 -1906
rect 1830 -2008 1864 -1974
rect 1830 -2076 1864 -2042
rect 1830 -2144 1864 -2110
rect 1830 -2212 1864 -2178
rect 1830 -2280 1864 -2246
rect 2894 -1396 2928 -1362
rect 2894 -1464 2928 -1430
rect 2894 -1532 2928 -1498
rect 2894 -1600 2928 -1566
rect 2894 -1668 2928 -1634
rect 2894 -1736 2928 -1702
rect 2894 -1804 2928 -1770
rect 2894 -1872 2928 -1838
rect 2894 -1940 2928 -1906
rect 2894 -2008 2928 -1974
rect 2894 -2076 2928 -2042
rect 2894 -2144 2928 -2110
rect 2894 -2212 2928 -2178
rect 2894 -2280 2928 -2246
rect 3958 -1396 3992 -1362
rect 3958 -1464 3992 -1430
rect 3958 -1532 3992 -1498
rect 3958 -1600 3992 -1566
rect 3958 -1668 3992 -1634
rect 3958 -1736 3992 -1702
rect 3958 -1804 3992 -1770
rect 3958 -1872 3992 -1838
rect 3958 -1940 3992 -1906
rect 3958 -2008 3992 -1974
rect 3958 -2076 3992 -2042
rect 3958 -2144 3992 -2110
rect 3958 -2212 3992 -2178
rect 3958 -2280 3992 -2246
rect -5266 -2410 -5232 -2376
rect -5266 -2478 -5232 -2444
rect -5266 -2546 -5232 -2512
rect -5266 -2614 -5232 -2580
rect -5266 -2682 -5232 -2648
<< locali >>
rect -3130 -1320 -3096 -1304
rect -5266 -1544 -5232 -1528
rect -4356 -1898 -4322 -1882
rect -3130 -2112 -3096 -2096
rect -2066 -1320 -2032 -1304
rect -2066 -2112 -2032 -2096
rect -1002 -1320 -968 -1304
rect -1002 -2112 -968 -2096
rect -298 -1320 -264 -1304
rect -298 -2312 -264 -2296
rect 766 -1320 800 -1304
rect 766 -2312 800 -2296
rect 1830 -1320 1864 -1304
rect 1830 -2312 1864 -2296
rect 2894 -1320 2928 -1304
rect 2894 -2312 2928 -2296
rect 3958 -1320 3992 -1304
rect 3958 -2312 3992 -2296
rect -5266 -2360 -5232 -2344
rect -5266 -2752 -5232 -2736
rect -3130 -2874 -3096 -2858
rect -5266 -2972 -5232 -2956
rect -5266 -3064 -5232 -3048
rect -3130 -3666 -3096 -3650
rect -2066 -2874 -2032 -2858
rect -2066 -3666 -2032 -3650
rect -1002 -2874 -968 -2858
rect 2 -2948 36 -2932
rect 2 -3140 36 -3126
rect 466 -2948 500 -2932
rect 466 -3140 500 -3126
rect 1530 -2948 1564 -2932
rect 1530 -3140 1564 -3126
rect 2130 -2948 2164 -2932
rect 2130 -3140 2164 -3126
rect 2594 -2948 2628 -2932
rect 2594 -3140 2628 -3126
rect 3658 -2948 3692 -2932
rect 3658 -3140 3692 -3126
rect -1002 -3666 -968 -3650
rect 1292 -3892 1326 -3876
rect -2766 -4414 -2762 -4198
rect -2766 -4482 -2760 -4414
rect -2480 -4482 -2474 -4198
rect -2766 -4488 -2474 -4482
rect -1572 -4482 -1566 -4474
rect -1290 -4482 -1284 -4474
rect -1572 -4488 -1284 -4482
rect 1292 -4884 1326 -4868
rect 2356 -3892 2390 -3876
rect 2356 -4884 2390 -4868
<< viali >>
rect -3130 -1366 -3096 -1320
rect -3130 -1400 -3096 -1366
rect -3130 -1434 -3096 -1400
rect -3130 -1468 -3096 -1434
rect -3130 -1502 -3096 -1468
rect -5266 -1560 -5232 -1544
rect -5266 -1594 -5232 -1560
rect -5266 -1628 -5232 -1594
rect -5266 -1662 -5232 -1628
rect -5266 -1696 -5232 -1662
rect -5266 -1730 -5232 -1696
rect -5266 -1764 -5232 -1730
rect -5266 -1798 -5232 -1764
rect -5266 -1832 -5232 -1798
rect -5266 -1866 -5232 -1832
rect -5266 -1920 -5232 -1866
rect -4356 -1560 -4322 -1506
rect -4356 -1594 -4322 -1560
rect -4356 -1628 -4322 -1594
rect -4356 -1662 -4322 -1628
rect -4356 -1696 -4322 -1662
rect -4356 -1730 -4322 -1696
rect -4356 -1764 -4322 -1730
rect -4356 -1798 -4322 -1764
rect -4356 -1832 -4322 -1798
rect -4356 -1866 -4322 -1832
rect -4356 -1882 -4322 -1866
rect -3130 -1536 -3096 -1502
rect -3130 -1570 -3096 -1536
rect -3130 -1604 -3096 -1570
rect -3130 -1638 -3096 -1604
rect -3130 -1672 -3096 -1638
rect -3130 -1706 -3096 -1672
rect -3130 -1740 -3096 -1706
rect -3130 -1774 -3096 -1740
rect -3130 -1808 -3096 -1774
rect -3130 -1842 -3096 -1808
rect -3130 -1876 -3096 -1842
rect -3130 -1910 -3096 -1876
rect -3130 -1944 -3096 -1910
rect -3130 -1978 -3096 -1944
rect -3130 -2012 -3096 -1978
rect -3130 -2046 -3096 -2012
rect -3130 -2080 -3096 -2046
rect -3130 -2096 -3096 -2080
rect -2066 -1366 -2032 -1320
rect -2066 -1400 -2032 -1366
rect -2066 -1434 -2032 -1400
rect -2066 -1468 -2032 -1434
rect -2066 -1502 -2032 -1468
rect -2066 -1536 -2032 -1502
rect -2066 -1570 -2032 -1536
rect -2066 -1604 -2032 -1570
rect -2066 -1638 -2032 -1604
rect -2066 -1672 -2032 -1638
rect -2066 -1706 -2032 -1672
rect -2066 -1740 -2032 -1706
rect -2066 -1774 -2032 -1740
rect -2066 -1808 -2032 -1774
rect -2066 -1842 -2032 -1808
rect -2066 -1876 -2032 -1842
rect -2066 -1910 -2032 -1876
rect -2066 -1944 -2032 -1910
rect -2066 -1978 -2032 -1944
rect -2066 -2012 -2032 -1978
rect -2066 -2046 -2032 -2012
rect -2066 -2080 -2032 -2046
rect -2066 -2096 -2032 -2080
rect -1002 -1366 -968 -1320
rect -1002 -1400 -968 -1366
rect -1002 -1434 -968 -1400
rect -1002 -1468 -968 -1434
rect -1002 -1502 -968 -1468
rect -1002 -1536 -968 -1502
rect -1002 -1570 -968 -1536
rect -1002 -1604 -968 -1570
rect -1002 -1638 -968 -1604
rect -1002 -1672 -968 -1638
rect -1002 -1706 -968 -1672
rect -1002 -1740 -968 -1706
rect -1002 -1774 -968 -1740
rect -1002 -1808 -968 -1774
rect -1002 -1842 -968 -1808
rect -1002 -1876 -968 -1842
rect -1002 -1910 -968 -1876
rect -1002 -1944 -968 -1910
rect -1002 -1978 -968 -1944
rect -1002 -2012 -968 -1978
rect -1002 -2046 -968 -2012
rect -1002 -2080 -968 -2046
rect -1002 -2096 -968 -2080
rect -298 -1362 -264 -1320
rect -298 -1396 -264 -1362
rect -298 -1430 -264 -1396
rect -298 -1464 -264 -1430
rect -298 -1498 -264 -1464
rect -298 -1532 -264 -1498
rect -298 -1566 -264 -1532
rect -298 -1600 -264 -1566
rect -298 -1634 -264 -1600
rect -298 -1668 -264 -1634
rect -298 -1702 -264 -1668
rect -298 -1736 -264 -1702
rect -298 -1770 -264 -1736
rect -298 -1804 -264 -1770
rect -298 -1838 -264 -1804
rect -298 -1872 -264 -1838
rect -298 -1906 -264 -1872
rect -298 -1940 -264 -1906
rect -298 -1974 -264 -1940
rect -298 -2008 -264 -1974
rect -298 -2042 -264 -2008
rect -298 -2076 -264 -2042
rect -298 -2110 -264 -2076
rect -298 -2144 -264 -2110
rect -298 -2178 -264 -2144
rect -298 -2212 -264 -2178
rect -298 -2246 -264 -2212
rect -298 -2280 -264 -2246
rect -298 -2296 -264 -2280
rect 766 -1362 800 -1320
rect 766 -1396 800 -1362
rect 766 -1430 800 -1396
rect 766 -1464 800 -1430
rect 766 -1498 800 -1464
rect 766 -1532 800 -1498
rect 766 -1566 800 -1532
rect 766 -1600 800 -1566
rect 766 -1634 800 -1600
rect 766 -1668 800 -1634
rect 766 -1702 800 -1668
rect 766 -1736 800 -1702
rect 766 -1770 800 -1736
rect 766 -1804 800 -1770
rect 766 -1838 800 -1804
rect 766 -1872 800 -1838
rect 766 -1906 800 -1872
rect 766 -1940 800 -1906
rect 766 -1974 800 -1940
rect 766 -2008 800 -1974
rect 766 -2042 800 -2008
rect 766 -2076 800 -2042
rect 766 -2110 800 -2076
rect 766 -2144 800 -2110
rect 766 -2178 800 -2144
rect 766 -2212 800 -2178
rect 766 -2246 800 -2212
rect 766 -2280 800 -2246
rect 766 -2296 800 -2280
rect 1830 -1362 1864 -1320
rect 1830 -1396 1864 -1362
rect 1830 -1430 1864 -1396
rect 1830 -1464 1864 -1430
rect 1830 -1498 1864 -1464
rect 1830 -1532 1864 -1498
rect 1830 -1566 1864 -1532
rect 1830 -1600 1864 -1566
rect 1830 -1634 1864 -1600
rect 1830 -1668 1864 -1634
rect 1830 -1702 1864 -1668
rect 1830 -1736 1864 -1702
rect 1830 -1770 1864 -1736
rect 1830 -1804 1864 -1770
rect 1830 -1838 1864 -1804
rect 1830 -1872 1864 -1838
rect 1830 -1906 1864 -1872
rect 1830 -1940 1864 -1906
rect 1830 -1974 1864 -1940
rect 1830 -2008 1864 -1974
rect 1830 -2042 1864 -2008
rect 1830 -2076 1864 -2042
rect 1830 -2110 1864 -2076
rect 1830 -2144 1864 -2110
rect 1830 -2178 1864 -2144
rect 1830 -2212 1864 -2178
rect 1830 -2246 1864 -2212
rect 1830 -2280 1864 -2246
rect 1830 -2296 1864 -2280
rect 2894 -1362 2928 -1320
rect 2894 -1396 2928 -1362
rect 2894 -1430 2928 -1396
rect 2894 -1464 2928 -1430
rect 2894 -1498 2928 -1464
rect 2894 -1532 2928 -1498
rect 2894 -1566 2928 -1532
rect 2894 -1600 2928 -1566
rect 2894 -1634 2928 -1600
rect 2894 -1668 2928 -1634
rect 2894 -1702 2928 -1668
rect 2894 -1736 2928 -1702
rect 2894 -1770 2928 -1736
rect 2894 -1804 2928 -1770
rect 2894 -1838 2928 -1804
rect 2894 -1872 2928 -1838
rect 2894 -1906 2928 -1872
rect 2894 -1940 2928 -1906
rect 2894 -1974 2928 -1940
rect 2894 -2008 2928 -1974
rect 2894 -2042 2928 -2008
rect 2894 -2076 2928 -2042
rect 2894 -2110 2928 -2076
rect 2894 -2144 2928 -2110
rect 2894 -2178 2928 -2144
rect 2894 -2212 2928 -2178
rect 2894 -2246 2928 -2212
rect 2894 -2280 2928 -2246
rect 2894 -2296 2928 -2280
rect 3958 -1362 3992 -1320
rect 3958 -1396 3992 -1362
rect 3958 -1430 3992 -1396
rect 3958 -1464 3992 -1430
rect 3958 -1498 3992 -1464
rect 3958 -1532 3992 -1498
rect 3958 -1566 3992 -1532
rect 3958 -1600 3992 -1566
rect 3958 -1634 3992 -1600
rect 3958 -1668 3992 -1634
rect 3958 -1702 3992 -1668
rect 3958 -1736 3992 -1702
rect 3958 -1770 3992 -1736
rect 3958 -1804 3992 -1770
rect 3958 -1838 3992 -1804
rect 3958 -1872 3992 -1838
rect 3958 -1906 3992 -1872
rect 3958 -1940 3992 -1906
rect 3958 -1974 3992 -1940
rect 3958 -2008 3992 -1974
rect 3958 -2042 3992 -2008
rect 3958 -2076 3992 -2042
rect 3958 -2110 3992 -2076
rect 3958 -2144 3992 -2110
rect 3958 -2178 3992 -2144
rect 3958 -2212 3992 -2178
rect 3958 -2246 3992 -2212
rect 3958 -2280 3992 -2246
rect 3958 -2296 3992 -2280
rect -5266 -2376 -5232 -2360
rect -5266 -2410 -5232 -2376
rect -5266 -2444 -5232 -2410
rect -5266 -2478 -5232 -2444
rect -5266 -2512 -5232 -2478
rect -5266 -2546 -5232 -2512
rect -5266 -2580 -5232 -2546
rect -5266 -2614 -5232 -2580
rect -5266 -2648 -5232 -2614
rect -5266 -2682 -5232 -2648
rect -5266 -2736 -5232 -2682
rect -3130 -2920 -3096 -2874
rect -3130 -2954 -3096 -2920
rect -5266 -2986 -5232 -2972
rect -5266 -3032 -5232 -2986
rect -5266 -3048 -5232 -3032
rect -3130 -2988 -3096 -2954
rect -3130 -3022 -3096 -2988
rect -3130 -3056 -3096 -3022
rect -3130 -3090 -3096 -3056
rect -3130 -3124 -3096 -3090
rect -3130 -3158 -3096 -3124
rect -3130 -3192 -3096 -3158
rect -3130 -3226 -3096 -3192
rect -3130 -3260 -3096 -3226
rect -3130 -3294 -3096 -3260
rect -3130 -3328 -3096 -3294
rect -3130 -3362 -3096 -3328
rect -3130 -3396 -3096 -3362
rect -3130 -3430 -3096 -3396
rect -3130 -3464 -3096 -3430
rect -3130 -3498 -3096 -3464
rect -3130 -3532 -3096 -3498
rect -3130 -3566 -3096 -3532
rect -3130 -3600 -3096 -3566
rect -3130 -3634 -3096 -3600
rect -3130 -3650 -3096 -3634
rect -2066 -2920 -2032 -2874
rect -2066 -2954 -2032 -2920
rect -2066 -2988 -2032 -2954
rect -2066 -3022 -2032 -2988
rect -2066 -3056 -2032 -3022
rect -2066 -3090 -2032 -3056
rect -2066 -3124 -2032 -3090
rect -2066 -3158 -2032 -3124
rect -2066 -3192 -2032 -3158
rect -2066 -3226 -2032 -3192
rect -2066 -3260 -2032 -3226
rect -2066 -3294 -2032 -3260
rect -2066 -3328 -2032 -3294
rect -2066 -3362 -2032 -3328
rect -2066 -3396 -2032 -3362
rect -2066 -3430 -2032 -3396
rect -2066 -3464 -2032 -3430
rect -2066 -3498 -2032 -3464
rect -2066 -3532 -2032 -3498
rect -2066 -3566 -2032 -3532
rect -2066 -3600 -2032 -3566
rect -2066 -3634 -2032 -3600
rect -2066 -3650 -2032 -3634
rect -1002 -2920 -968 -2874
rect -1002 -2954 -968 -2920
rect -1002 -2988 -968 -2954
rect -1002 -3022 -968 -2988
rect -1002 -3056 -968 -3022
rect -1002 -3090 -968 -3056
rect -1002 -3124 -968 -3090
rect -1002 -3158 -968 -3124
rect 2 -2990 36 -2948
rect 2 -3024 36 -2990
rect 2 -3058 36 -3024
rect 2 -3092 36 -3058
rect 2 -3126 36 -3092
rect 466 -2990 500 -2948
rect 466 -3024 500 -2990
rect 466 -3058 500 -3024
rect 466 -3092 500 -3058
rect 466 -3126 500 -3092
rect 1530 -2990 1564 -2948
rect 1530 -3024 1564 -2990
rect 1530 -3058 1564 -3024
rect 1530 -3092 1564 -3058
rect 1530 -3126 1564 -3092
rect 2130 -2990 2164 -2948
rect 2130 -3024 2164 -2990
rect 2130 -3058 2164 -3024
rect 2130 -3092 2164 -3058
rect 2130 -3126 2164 -3092
rect 2594 -2990 2628 -2948
rect 2594 -3024 2628 -2990
rect 2594 -3058 2628 -3024
rect 2594 -3092 2628 -3058
rect 2594 -3126 2628 -3092
rect 3658 -2990 3692 -2948
rect 3658 -3024 3692 -2990
rect 3658 -3058 3692 -3024
rect 3658 -3092 3692 -3058
rect 3658 -3126 3692 -3092
rect -1002 -3192 -968 -3158
rect -1002 -3226 -968 -3192
rect -1002 -3260 -968 -3226
rect -1002 -3294 -968 -3260
rect -1002 -3328 -968 -3294
rect -1002 -3362 -968 -3328
rect -1002 -3396 -968 -3362
rect -1002 -3430 -968 -3396
rect -1002 -3464 -968 -3430
rect -1002 -3498 -968 -3464
rect -1002 -3532 -968 -3498
rect -1002 -3566 -968 -3532
rect -1002 -3600 -968 -3566
rect -1002 -3634 -968 -3600
rect -1002 -3650 -968 -3634
rect 1292 -3934 1326 -3892
rect 1292 -3968 1326 -3934
rect -2972 -4048 -2270 -3988
rect -2972 -4632 -2910 -4048
rect -2824 -4198 -2416 -4138
rect -2824 -4488 -2766 -4198
rect -2474 -4488 -2416 -4198
rect -2824 -4542 -2416 -4488
rect -2332 -4632 -2270 -4048
rect -2972 -4692 -2270 -4632
rect -1778 -4048 -1076 -3988
rect -1778 -4632 -1716 -4048
rect -1630 -4198 -1222 -4138
rect -1630 -4488 -1572 -4198
rect -1284 -4488 -1222 -4198
rect -1630 -4542 -1222 -4488
rect -1138 -4632 -1076 -4048
rect -1778 -4692 -1076 -4632
rect 1292 -4002 1326 -3968
rect 1292 -4036 1326 -4002
rect 1292 -4070 1326 -4036
rect 1292 -4104 1326 -4070
rect 1292 -4138 1326 -4104
rect 1292 -4172 1326 -4138
rect 1292 -4206 1326 -4172
rect 1292 -4240 1326 -4206
rect 1292 -4274 1326 -4240
rect 1292 -4308 1326 -4274
rect 1292 -4342 1326 -4308
rect 1292 -4376 1326 -4342
rect 1292 -4410 1326 -4376
rect 1292 -4444 1326 -4410
rect 1292 -4478 1326 -4444
rect 1292 -4512 1326 -4478
rect 1292 -4546 1326 -4512
rect 1292 -4580 1326 -4546
rect 1292 -4614 1326 -4580
rect 1292 -4648 1326 -4614
rect 1292 -4682 1326 -4648
rect 1292 -4716 1326 -4682
rect 1292 -4750 1326 -4716
rect 1292 -4784 1326 -4750
rect 1292 -4818 1326 -4784
rect 1292 -4852 1326 -4818
rect 1292 -4868 1326 -4852
rect 2356 -3934 2390 -3892
rect 2356 -3968 2390 -3934
rect 2356 -4002 2390 -3968
rect 2356 -4036 2390 -4002
rect 2356 -4070 2390 -4036
rect 2356 -4104 2390 -4070
rect 2356 -4138 2390 -4104
rect 2356 -4172 2390 -4138
rect 2356 -4206 2390 -4172
rect 2356 -4240 2390 -4206
rect 2356 -4274 2390 -4240
rect 2356 -4308 2390 -4274
rect 2356 -4342 2390 -4308
rect 2356 -4376 2390 -4342
rect 2356 -4410 2390 -4376
rect 2356 -4444 2390 -4410
rect 2356 -4478 2390 -4444
rect 2356 -4512 2390 -4478
rect 2356 -4546 2390 -4512
rect 2356 -4580 2390 -4546
rect 2356 -4614 2390 -4580
rect 2356 -4648 2390 -4614
rect 2356 -4682 2390 -4648
rect 2356 -4716 2390 -4682
rect 2356 -4750 2390 -4716
rect 2356 -4784 2390 -4750
rect 2356 -4818 2390 -4784
rect 2356 -4852 2390 -4818
rect 2356 -4868 2390 -4852
<< metal1 >>
rect -5328 52 -5170 58
rect -5748 -1494 -5742 -1442
rect -5374 -1494 -5368 -1442
rect -5328 -1526 -5170 -398
rect -4362 52 -4242 58
rect -5136 -1494 -5130 -1442
rect -4762 -1494 -4668 -1442
rect -5328 -1528 -5152 -1526
rect -5830 -2748 -5776 -1532
rect -5346 -1544 -5152 -1528
rect -4734 -1532 -4668 -1494
rect -5346 -1920 -5266 -1544
rect -5232 -1920 -5152 -1544
rect -5346 -1932 -5152 -1920
rect -5742 -2310 -5736 -2258
rect -5368 -2310 -5362 -2258
rect -5354 -2882 -5300 -2348
rect -5272 -2360 -5226 -1932
rect -5272 -2736 -5266 -2360
rect -5232 -2736 -5226 -2360
rect -5272 -2748 -5226 -2736
rect -5198 -2310 -5192 -2258
rect -4762 -2310 -4756 -2258
rect -5386 -2928 -5300 -2882
rect -5812 -5314 -5758 -2960
rect -5354 -3060 -5300 -2928
rect -5198 -2882 -5144 -2310
rect -4722 -2748 -4668 -1532
rect -4362 -1506 -4242 -398
rect -304 52 -184 58
rect -3672 -1320 -3616 -1308
rect -3224 -1320 -3172 -1314
rect -3136 -1320 -3090 -1308
rect -3054 -1318 -3002 -1312
rect -4362 -1882 -4356 -1506
rect -4322 -1882 -4242 -1506
rect -4362 -1894 -4242 -1882
rect -3830 -1506 -3778 -1500
rect -3830 -1888 -3778 -1882
rect -4274 -1984 -4220 -1932
rect -3852 -1984 -3846 -1932
rect -4274 -2258 -4222 -1984
rect -3672 -2072 -3670 -1320
rect -3618 -2072 -3616 -1320
rect -3672 -2138 -3616 -2072
rect -3226 -2096 -3224 -1320
rect -3172 -2096 -3170 -1320
rect -3226 -2106 -3170 -2096
rect -3136 -2096 -3130 -1320
rect -3096 -2096 -3090 -1320
rect -3680 -2190 -3674 -2138
rect -3232 -2190 -3226 -2138
rect -4280 -2310 -4274 -2258
rect -4222 -2310 -4216 -2258
rect -3136 -2874 -3090 -2096
rect -3056 -2096 -3054 -1318
rect -3002 -2096 -3000 -1318
rect -3056 -2102 -3000 -2096
rect -2606 -1320 -2554 -1314
rect -2606 -2102 -2554 -2096
rect -2162 -1318 -2106 -1312
rect -2162 -2090 -2160 -1318
rect -2108 -2090 -2106 -1318
rect -2162 -2100 -2106 -2090
rect -2072 -1320 -2026 -1308
rect -2072 -2096 -2066 -1320
rect -2032 -2096 -2026 -1320
rect -3000 -2190 -2994 -2138
rect -2626 -2190 -2620 -2138
rect -2542 -2190 -2536 -2138
rect -2168 -2190 -2162 -2138
rect -3000 -2780 -2626 -2190
rect -2536 -2780 -2162 -2190
rect -3000 -2832 -2994 -2780
rect -2626 -2832 -2620 -2780
rect -2542 -2832 -2536 -2780
rect -2168 -2832 -2162 -2780
rect -5198 -2928 -5124 -2882
rect -5266 -2960 -5232 -2956
rect -5272 -2972 -5226 -2960
rect -5272 -3048 -5266 -2972
rect -5232 -3048 -5226 -2972
rect -5272 -5308 -5226 -3048
rect -5198 -3754 -5144 -2928
rect -5198 -3852 -5144 -3846
rect -5812 -5770 -5758 -5764
rect -5276 -5314 -5222 -5308
rect -5276 -5770 -5222 -5764
rect -4748 -5314 -4694 -2960
rect -4748 -5770 -4694 -5764
rect -3136 -3650 -3130 -2874
rect -3096 -3650 -3090 -2874
rect -3136 -5308 -3090 -3650
rect -3056 -2874 -3000 -2864
rect -3056 -3650 -3054 -2874
rect -3002 -3650 -3000 -2874
rect -3056 -3656 -3000 -3650
rect -2606 -2874 -2554 -2868
rect -2162 -2874 -2106 -2864
rect -2162 -3646 -2160 -2874
rect -2108 -3646 -2106 -2874
rect -2072 -2874 -2026 -2096
rect -1992 -1318 -1936 -1312
rect -1992 -2096 -1990 -1318
rect -1938 -2096 -1936 -1318
rect -1992 -2106 -1936 -2096
rect -1542 -1320 -1490 -1314
rect -1542 -2102 -1490 -2096
rect -1098 -1318 -1042 -1312
rect -1098 -2090 -1096 -1318
rect -1044 -2090 -1042 -1318
rect -1098 -2100 -1042 -2090
rect -1008 -1320 -962 -1308
rect -1008 -2096 -1002 -1320
rect -968 -2096 -962 -1320
rect -1936 -2190 -1930 -2138
rect -1562 -2190 -1556 -2138
rect -1478 -2190 -1472 -2138
rect -1104 -2190 -1098 -2138
rect -1936 -2780 -1562 -2190
rect -1472 -2780 -1098 -2190
rect -1936 -2832 -1930 -2780
rect -1562 -2832 -1556 -2780
rect -1478 -2832 -1472 -2780
rect -1104 -2832 -1098 -2780
rect -2606 -3656 -2554 -3650
rect -2160 -3652 -2108 -3646
rect -2072 -3650 -2066 -2874
rect -2032 -3650 -2026 -2874
rect -1992 -2874 -1936 -2864
rect -1992 -3646 -1990 -2874
rect -1938 -3646 -1936 -2874
rect -1542 -2874 -1490 -2868
rect -2984 -3988 -2258 -3982
rect -2984 -4692 -2972 -3988
rect -2910 -4138 -2332 -4048
rect -2910 -4542 -2824 -4138
rect -2766 -4204 -2474 -4198
rect -2766 -4482 -2760 -4204
rect -2692 -4274 -2548 -4268
rect -2692 -4406 -2686 -4274
rect -2554 -4406 -2548 -4274
rect -2692 -4412 -2548 -4406
rect -2480 -4482 -2474 -4204
rect -2766 -4488 -2474 -4482
rect -2416 -4542 -2332 -4138
rect -2910 -4632 -2332 -4542
rect -2270 -4692 -2258 -3988
rect -3136 -5314 -3084 -5308
rect -3136 -5770 -3084 -5764
rect -2984 -5314 -2258 -4692
rect -2984 -5770 -2258 -5764
rect -2072 -5308 -2026 -3650
rect -1990 -3652 -1938 -3646
rect -1098 -2874 -1042 -2864
rect -1098 -3650 -1096 -2874
rect -1044 -3650 -1042 -2874
rect -1008 -2874 -962 -2096
rect -928 -1318 -872 -1312
rect -928 -2096 -926 -1318
rect -874 -2096 -872 -1318
rect -928 -2106 -872 -2096
rect -478 -1320 -426 -1314
rect -478 -2102 -426 -2096
rect -304 -1320 -184 -398
rect 722 52 842 58
rect -872 -2190 -866 -2138
rect -498 -2190 -492 -2138
rect -872 -2780 -498 -2190
rect -304 -2296 -298 -1320
rect -264 -2296 -184 -1320
rect -304 -2308 -184 -2296
rect 224 -1320 276 -1314
rect 224 -2302 276 -2296
rect 722 -1320 842 -398
rect 1786 52 1906 58
rect 722 -2296 766 -1320
rect 800 -2296 842 -1320
rect 722 -2308 842 -2296
rect 1286 -2346 1344 -1308
rect 1786 -1320 1906 -398
rect 2850 52 2970 58
rect 1786 -2296 1830 -1320
rect 1864 -2296 1906 -1320
rect 1786 -2308 1906 -2296
rect 2350 -1320 2406 -1310
rect 2350 -2296 2352 -1320
rect 2404 -2296 2406 -1320
rect 2350 -2306 2406 -2296
rect 2850 -1320 2970 -398
rect 3878 52 3998 58
rect 2850 -2296 2894 -1320
rect 2928 -2296 2970 -1320
rect 2850 -2308 2970 -2296
rect 3414 -2346 3472 -1308
rect 3878 -1320 3998 -398
rect 3878 -2296 3958 -1320
rect 3992 -2296 3998 -1320
rect 3878 -2308 3998 -2296
rect -184 -2398 -178 -2346
rect 3916 -2398 3922 -2346
rect 126 -2534 132 -2430
rect 364 -2534 370 -2430
rect 2254 -2534 2260 -2430
rect 2492 -2534 2498 -2430
rect -230 -2678 -224 -2574
rect -120 -2678 -114 -2574
rect -224 -2718 -120 -2678
rect -872 -2832 -866 -2780
rect -498 -2832 -492 -2780
rect -230 -2822 -224 -2718
rect -120 -2822 -114 -2718
rect 132 -2854 370 -2534
rect 590 -2822 596 -2718
rect 1428 -2822 1434 -2718
rect -1008 -3650 -1002 -2874
rect -968 -3650 -962 -2874
rect -928 -2874 -872 -2864
rect -928 -3648 -926 -2874
rect -874 -3648 -872 -2874
rect -478 -2874 -426 -2868
rect -1542 -3656 -1490 -3650
rect -1096 -3656 -1044 -3650
rect -1790 -3988 -1064 -3982
rect -1790 -4692 -1778 -3988
rect -1716 -4138 -1138 -4048
rect -1716 -4542 -1630 -4138
rect -1572 -4204 -1284 -4198
rect -1572 -4482 -1566 -4204
rect -1498 -4274 -1354 -4268
rect -1498 -4406 -1492 -4274
rect -1360 -4406 -1354 -4274
rect -1498 -4412 -1354 -4406
rect -1290 -4482 -1284 -4204
rect -1572 -4488 -1284 -4482
rect -1222 -4542 -1138 -4138
rect -1716 -4632 -1138 -4542
rect -1076 -4692 -1064 -3988
rect -2072 -5314 -2020 -5308
rect -2072 -5770 -2020 -5764
rect -1790 -5314 -1064 -4692
rect -1790 -5770 -1064 -5764
rect -1008 -5308 -962 -3650
rect -926 -3654 -874 -3648
rect 132 -2906 138 -2854
rect 206 -2864 296 -2854
rect 206 -2906 212 -2864
rect 290 -2906 296 -2864
rect 364 -2906 370 -2854
rect 596 -2854 1434 -2822
rect 596 -2906 602 -2854
rect 970 -2866 1060 -2854
rect 970 -2906 976 -2866
rect 1054 -2906 1060 -2866
rect 1428 -2906 1434 -2854
rect 2260 -2854 2498 -2534
rect 4168 -2678 4174 -2574
rect 4336 -2678 4348 -2574
rect 2718 -2822 2724 -2718
rect 3556 -2822 3562 -2718
rect 2730 -2854 3556 -2822
rect 2260 -2906 2266 -2854
rect 2334 -2860 2424 -2854
rect 2334 -2906 2340 -2860
rect 2418 -2906 2424 -2860
rect 2492 -2906 2498 -2854
rect 2724 -2906 2730 -2854
rect 3098 -2866 3188 -2854
rect 3098 -2906 3104 -2866
rect 3182 -2906 3188 -2866
rect 3556 -2906 3562 -2854
rect -478 -3656 -426 -3650
rect -4 -2948 42 -2936
rect -4 -3126 2 -2948
rect 36 -3126 42 -2948
rect -4 -3604 42 -3126
rect 70 -3458 126 -2936
rect 222 -2948 278 -2938
rect 276 -3136 278 -2948
rect 222 -3142 278 -3136
rect 376 -3458 432 -2936
rect 70 -3562 76 -3458
rect 128 -3562 134 -3458
rect 368 -3562 374 -3458
rect 426 -3562 432 -3458
rect 460 -2948 506 -2936
rect 460 -3126 466 -2948
rect 500 -3126 506 -2948
rect 460 -3604 506 -3126
rect 534 -3458 590 -2936
rect 986 -2948 1042 -2938
rect 986 -3136 988 -2948
rect 1040 -3136 1042 -2948
rect 988 -3142 1040 -3136
rect 1440 -3458 1496 -2936
rect 534 -3562 540 -3458
rect 592 -3562 598 -3458
rect 722 -3562 728 -3458
rect 780 -3562 786 -3458
rect 1432 -3562 1438 -3458
rect 1490 -3562 1496 -3458
rect 1524 -2948 1570 -2936
rect 1524 -3126 1530 -2948
rect 1564 -3126 1570 -2948
rect -4 -3708 2 -3604
rect 54 -3708 60 -3604
rect 452 -3708 458 -3604
rect 510 -3708 516 -3604
rect 726 -3880 782 -3562
rect 1524 -3604 1570 -3126
rect 2124 -2948 2170 -2936
rect 2124 -3126 2130 -2948
rect 2164 -3126 2170 -2948
rect 2124 -3604 2170 -3126
rect 2198 -3458 2254 -2936
rect 2350 -2948 2406 -2938
rect 2404 -3136 2406 -2948
rect 2350 -3142 2404 -3136
rect 2504 -3458 2560 -2936
rect 2198 -3562 2204 -3458
rect 2256 -3562 2262 -3458
rect 2496 -3562 2502 -3458
rect 2554 -3562 2560 -3458
rect 2588 -2948 2634 -2936
rect 2588 -3126 2594 -2948
rect 2628 -3126 2634 -2948
rect 2588 -3604 2634 -3126
rect 2662 -3458 2718 -2936
rect 3114 -2948 3170 -2938
rect 3114 -3136 3116 -2948
rect 3168 -3136 3170 -2948
rect 3116 -3142 3168 -3136
rect 3568 -3458 3624 -2936
rect 2662 -3562 2668 -3458
rect 2720 -3562 2726 -3458
rect 2896 -3562 2902 -3458
rect 2954 -3562 2960 -3458
rect 3560 -3562 3566 -3458
rect 3618 -3562 3624 -3458
rect 3652 -2948 3698 -2936
rect 3652 -3126 3658 -2948
rect 3692 -3126 3698 -2948
rect 1278 -3708 1284 -3604
rect 1336 -3708 1342 -3604
rect 1516 -3708 1522 -3604
rect 1574 -3708 1580 -3604
rect 2116 -3708 2122 -3604
rect 2174 -3708 2180 -3604
rect 2342 -3708 2348 -3604
rect 2400 -3708 2406 -3604
rect 2580 -3708 2586 -3604
rect 2638 -3708 2644 -3604
rect 816 -3852 822 -3800
rect 1190 -3852 1196 -3800
rect 1286 -3880 1332 -3708
rect 1422 -3852 1428 -3800
rect 1796 -3852 1802 -3800
rect 1880 -3852 1886 -3800
rect 2254 -3852 2260 -3800
rect 2350 -3880 2396 -3708
rect 2486 -3852 2492 -3800
rect 2860 -3852 2866 -3800
rect 2900 -3880 2956 -3562
rect 3652 -3604 3698 -3126
rect 3634 -3708 3640 -3604
rect 3692 -3708 3698 -3604
rect 726 -4880 800 -3880
rect 1212 -3892 1406 -3880
rect 1212 -4868 1292 -3892
rect 1326 -4868 1406 -3892
rect 1212 -4880 1406 -4868
rect 1812 -3890 1868 -3880
rect 1812 -4866 1814 -3890
rect 1866 -4866 1868 -3890
rect 1812 -4876 1868 -4866
rect 2276 -3892 2470 -3880
rect 2276 -4868 2356 -3892
rect 2390 -4868 2470 -3892
rect 2276 -4880 2470 -4868
rect 2882 -4880 2956 -3880
rect 4174 -4880 4348 -2678
rect -1008 -5314 -956 -5308
rect -1008 -5770 -956 -5764
rect 1248 -5314 1368 -4880
rect 1248 -5770 1368 -5764
rect 2312 -5314 2432 -4880
rect 2312 -5770 2432 -5764
<< via1 >>
rect -5328 -398 -5170 52
rect -5742 -1494 -5374 -1442
rect -4362 -398 -4242 52
rect -5130 -1494 -4762 -1442
rect -5736 -2310 -5368 -2258
rect -5192 -2310 -4762 -2258
rect -304 -398 -184 52
rect -3830 -1882 -3778 -1506
rect -4220 -1984 -3852 -1932
rect -3670 -2072 -3618 -1320
rect -3224 -2096 -3172 -1320
rect -3674 -2190 -3232 -2138
rect -4274 -2310 -4222 -2258
rect -3054 -2096 -3002 -1318
rect -2606 -2096 -2554 -1320
rect -2160 -2090 -2108 -1318
rect -2994 -2190 -2626 -2138
rect -2536 -2190 -2168 -2138
rect -2994 -2832 -2626 -2780
rect -2536 -2832 -2168 -2780
rect -5198 -3846 -5144 -3754
rect -5812 -5764 -5758 -5314
rect -5276 -5764 -5222 -5314
rect -4748 -5764 -4694 -5314
rect -3054 -3650 -3002 -2874
rect -2606 -3650 -2554 -2874
rect -2160 -3646 -2108 -2874
rect -1990 -2096 -1938 -1318
rect -1542 -2096 -1490 -1320
rect -1096 -2090 -1044 -1318
rect -1930 -2190 -1562 -2138
rect -1472 -2190 -1104 -2138
rect -1930 -2832 -1562 -2780
rect -1472 -2832 -1104 -2780
rect -1990 -3646 -1938 -2874
rect -2686 -4406 -2554 -4274
rect -3136 -5764 -3084 -5314
rect -2984 -5764 -2258 -5314
rect -1542 -3650 -1490 -2874
rect -1096 -3650 -1044 -2874
rect -926 -2096 -874 -1318
rect -478 -2096 -426 -1320
rect 722 -398 842 52
rect -866 -2190 -498 -2138
rect 224 -2296 276 -1320
rect 1786 -398 1906 52
rect 2850 -398 2970 52
rect 2352 -2296 2404 -1320
rect 3878 -398 3998 52
rect -178 -2398 3916 -2346
rect 132 -2534 364 -2430
rect 2260 -2534 2492 -2430
rect -224 -2678 -120 -2574
rect -866 -2832 -498 -2780
rect -224 -2822 -120 -2718
rect 596 -2822 1428 -2718
rect -926 -3648 -874 -2874
rect -1492 -4406 -1360 -4274
rect -2072 -5764 -2020 -5314
rect -1790 -5764 -1064 -5314
rect -478 -3650 -426 -2874
rect 138 -2906 206 -2854
rect 296 -2906 364 -2854
rect 602 -2906 970 -2854
rect 1060 -2906 1428 -2854
rect 4174 -2678 4336 -2574
rect 2724 -2822 3556 -2718
rect 2266 -2906 2334 -2854
rect 2424 -2906 2492 -2854
rect 2730 -2906 3098 -2854
rect 3188 -2906 3556 -2854
rect 222 -3136 276 -2948
rect 76 -3562 128 -3458
rect 374 -3562 426 -3458
rect 988 -3136 1040 -2948
rect 540 -3562 592 -3458
rect 728 -3562 780 -3458
rect 1438 -3562 1490 -3458
rect 2 -3708 54 -3604
rect 458 -3708 510 -3604
rect 2350 -3136 2404 -2948
rect 2204 -3562 2256 -3458
rect 2502 -3562 2554 -3458
rect 3116 -3136 3168 -2948
rect 2668 -3562 2720 -3458
rect 2902 -3562 2954 -3458
rect 3566 -3562 3618 -3458
rect 1284 -3708 1336 -3604
rect 1522 -3708 1574 -3604
rect 2122 -3708 2174 -3604
rect 2348 -3708 2400 -3604
rect 2586 -3708 2638 -3604
rect 822 -3852 1190 -3800
rect 1428 -3852 1796 -3800
rect 1886 -3852 2254 -3800
rect 2492 -3852 2860 -3800
rect 3640 -3708 3692 -3604
rect 1814 -4866 1866 -3890
rect -1008 -5764 -956 -5314
rect 1248 -5764 1368 -5314
rect 2312 -5764 2432 -5314
<< metal2 >>
rect -5848 52 4348 64
rect -5848 -398 -5328 52
rect -5170 -398 -4362 52
rect -4242 48 -304 52
rect -4242 -394 -2608 48
rect -2552 -394 -1544 48
rect -1488 -394 -480 48
rect -424 -394 -304 48
rect -4242 -398 -304 -394
rect -184 -398 722 52
rect 842 -398 1786 52
rect 1906 -398 2850 52
rect 2970 -398 3878 52
rect 3998 -398 4348 52
rect -5848 -404 4348 -398
rect -3670 -1320 -3618 -1314
rect -5748 -1494 -5742 -1442
rect -5374 -1494 -5130 -1442
rect -4762 -1494 -4756 -1442
rect -3830 -1506 -3670 -1500
rect -3778 -1882 -3670 -1506
rect -3830 -1894 -3670 -1882
rect -4226 -1984 -4220 -1932
rect -3852 -1984 -3846 -1932
rect -3670 -2078 -3618 -2072
rect -3226 -1320 -3170 -1310
rect -3226 -2106 -3170 -2096
rect -3056 -1318 -3000 -1308
rect -3056 -2106 -3000 -2096
rect -2608 -1320 -2552 -1310
rect -2608 -2106 -2552 -2096
rect -2162 -1318 -2106 -1308
rect -2162 -2100 -2106 -2090
rect -1992 -1318 -1936 -1308
rect -1992 -2106 -1936 -2096
rect -1544 -1320 -1488 -1310
rect -1544 -2106 -1488 -2096
rect -1098 -1318 -1042 -1308
rect -1098 -2100 -1042 -2090
rect -928 -1318 -872 -1308
rect -928 -2106 -872 -2096
rect -480 -1320 -424 -1310
rect -480 -2106 -424 -2096
rect 222 -1320 278 -1310
rect -3680 -2138 -486 -2134
rect -3680 -2190 -3674 -2138
rect -3232 -2190 -2994 -2138
rect -2626 -2190 -2536 -2138
rect -2168 -2190 -1930 -2138
rect -1562 -2190 -1472 -2138
rect -1104 -2190 -866 -2138
rect -498 -2190 -486 -2138
rect -3680 -2194 -486 -2190
rect -5742 -2310 -5736 -2258
rect -5368 -2310 -5192 -2258
rect -4762 -2310 -4274 -2258
rect -4222 -2310 -4216 -2258
rect 222 -2306 278 -2296
rect 2350 -1320 2406 -1310
rect 2350 -2306 2406 -2296
rect -184 -2344 3112 -2342
rect -184 -2346 984 -2344
rect 1044 -2346 3112 -2344
rect 3172 -2346 3922 -2342
rect -184 -2398 -178 -2346
rect 3916 -2398 3922 -2346
rect -184 -2400 984 -2398
rect 1044 -2400 3922 -2398
rect -184 -2402 3922 -2400
rect -3066 -2436 132 -2430
rect -3066 -2528 -3056 -2436
rect -3000 -2528 -2162 -2436
rect -2106 -2528 -1992 -2436
rect -1936 -2528 -1098 -2436
rect -1042 -2528 -928 -2436
rect -872 -2528 132 -2436
rect -3066 -2534 132 -2528
rect 364 -2534 2260 -2430
rect 2492 -2534 2498 -2430
rect -3236 -2580 -224 -2574
rect -3236 -2672 -3226 -2580
rect -3170 -2672 -224 -2580
rect -3236 -2678 -224 -2672
rect -120 -2678 -114 -2574
rect 212 -2580 4174 -2574
rect 212 -2672 222 -2580
rect 278 -2672 2350 -2580
rect 2406 -2672 4174 -2580
rect 212 -2678 4174 -2672
rect 4336 -2678 4342 -2574
rect -3006 -2780 -486 -2776
rect -3006 -2832 -2994 -2780
rect -2626 -2832 -2536 -2780
rect -2168 -2832 -1930 -2780
rect -1562 -2832 -1472 -2780
rect -1104 -2832 -866 -2780
rect -498 -2832 -486 -2780
rect -230 -2822 -224 -2718
rect -120 -2822 596 -2718
rect 1428 -2822 2724 -2718
rect 3556 -2822 3562 -2718
rect -3006 -2836 -486 -2832
rect 132 -2854 370 -2850
rect -3056 -2874 -3000 -2864
rect -3056 -3660 -3000 -3650
rect -2608 -2874 -2552 -2864
rect -2608 -3660 -2552 -3650
rect -2162 -2874 -2106 -2864
rect -2162 -3656 -2106 -3646
rect -1992 -2874 -1936 -2864
rect -1992 -3656 -1936 -3646
rect -1544 -2874 -1488 -2864
rect -1544 -3660 -1488 -3650
rect -1098 -2874 -1042 -2864
rect -1098 -3660 -1042 -3650
rect -928 -2874 -872 -2864
rect -928 -3658 -872 -3648
rect -480 -2874 -424 -2864
rect 132 -2906 138 -2854
rect 206 -2906 296 -2854
rect 364 -2906 370 -2854
rect 132 -2910 370 -2906
rect 596 -2854 1434 -2850
rect 596 -2906 602 -2854
rect 970 -2906 1060 -2854
rect 1428 -2906 1434 -2854
rect 596 -2910 1434 -2906
rect 2260 -2854 2498 -2850
rect 2260 -2906 2266 -2854
rect 2334 -2906 2424 -2854
rect 2492 -2906 2498 -2854
rect 2260 -2910 2498 -2906
rect 2724 -2854 3562 -2850
rect 2724 -2906 2730 -2854
rect 3098 -2906 3188 -2854
rect 3556 -2906 3562 -2854
rect 2724 -2910 3562 -2906
rect 222 -2948 278 -2938
rect 222 -3146 278 -3136
rect 986 -2948 1042 -2938
rect 986 -3146 1042 -3136
rect 2350 -2948 2406 -2938
rect 2350 -3146 2406 -3136
rect 3114 -2948 3170 -2938
rect 3114 -3146 3170 -3136
rect 70 -3562 76 -3458
rect 128 -3562 374 -3458
rect 426 -3562 540 -3458
rect 592 -3562 728 -3458
rect 780 -3562 1438 -3458
rect 1490 -3464 2204 -3458
rect 1490 -3556 1812 -3464
rect 1868 -3556 2204 -3464
rect 1490 -3562 2204 -3556
rect 2256 -3562 2502 -3458
rect 2554 -3562 2668 -3458
rect 2720 -3562 2902 -3458
rect 2954 -3562 3566 -3458
rect 3618 -3562 3624 -3458
rect -480 -3660 -424 -3650
rect -4 -3708 2 -3604
rect 54 -3708 458 -3604
rect 510 -3708 1284 -3604
rect 1336 -3708 1522 -3604
rect 1574 -3708 2122 -3604
rect 2174 -3708 2348 -3604
rect 2400 -3708 2586 -3604
rect 2638 -3708 3640 -3604
rect 3692 -3708 3698 -3604
rect -5198 -3754 2866 -3748
rect -5144 -3800 2866 -3754
rect -5144 -3846 822 -3800
rect -5198 -3852 822 -3846
rect 1190 -3852 1428 -3800
rect 1796 -3852 1886 -3800
rect 2254 -3852 2492 -3800
rect 2860 -3852 2866 -3800
rect 1812 -3890 1868 -3880
rect -2692 -4274 -2548 -4268
rect -1498 -4274 -1354 -4268
rect -3232 -4284 -2686 -4274
rect -3232 -4396 -3222 -4284
rect -3166 -4396 -2686 -4284
rect -3232 -4406 -2686 -4396
rect -2554 -4406 -2548 -4274
rect -1998 -4284 -1492 -4274
rect -1998 -4396 -1988 -4284
rect -1932 -4396 -1492 -4284
rect -1998 -4406 -1492 -4396
rect -1360 -4406 -1354 -4274
rect -2692 -4412 -2548 -4406
rect -1498 -4412 -1354 -4406
rect 1812 -4876 1868 -4866
rect -5848 -5314 4348 -5308
rect -5848 -5764 -5812 -5314
rect -5758 -5764 -5276 -5314
rect -5222 -5764 -4748 -5314
rect -4694 -5764 -3136 -5314
rect -3084 -5764 -2984 -5314
rect -2258 -5764 -2072 -5314
rect -2020 -5764 -1790 -5314
rect -1064 -5764 -1008 -5314
rect -956 -5764 1248 -5314
rect 1368 -5764 2312 -5314
rect 2432 -5764 4348 -5314
rect -5848 -5776 4348 -5764
<< via2 >>
rect -2608 -394 -2552 48
rect -1544 -394 -1488 48
rect -480 -394 -424 48
rect -3226 -2096 -3224 -1320
rect -3224 -2096 -3172 -1320
rect -3172 -2096 -3170 -1320
rect -3056 -2096 -3054 -1318
rect -3054 -2096 -3002 -1318
rect -3002 -2096 -3000 -1318
rect -2608 -2096 -2606 -1320
rect -2606 -2096 -2554 -1320
rect -2554 -2096 -2552 -1320
rect -2162 -2090 -2160 -1318
rect -2160 -2090 -2108 -1318
rect -2108 -2090 -2106 -1318
rect -1992 -2096 -1990 -1318
rect -1990 -2096 -1938 -1318
rect -1938 -2096 -1936 -1318
rect -1544 -2096 -1542 -1320
rect -1542 -2096 -1490 -1320
rect -1490 -2096 -1488 -1320
rect -1098 -2090 -1096 -1318
rect -1096 -2090 -1044 -1318
rect -1044 -2090 -1042 -1318
rect -928 -2096 -926 -1318
rect -926 -2096 -874 -1318
rect -874 -2096 -872 -1318
rect -480 -2096 -478 -1320
rect -478 -2096 -426 -1320
rect -426 -2096 -424 -1320
rect 222 -2296 224 -1320
rect 224 -2296 276 -1320
rect 276 -2296 278 -1320
rect 2350 -2296 2352 -1320
rect 2352 -2296 2404 -1320
rect 2404 -2296 2406 -1320
rect 984 -2346 1044 -2344
rect 3112 -2346 3172 -2342
rect 984 -2398 1044 -2346
rect 3112 -2398 3172 -2346
rect 984 -2400 1044 -2398
rect -3056 -2528 -3000 -2436
rect -2162 -2528 -2106 -2436
rect -1992 -2528 -1936 -2436
rect -1098 -2528 -1042 -2436
rect -928 -2528 -872 -2436
rect -3226 -2672 -3170 -2580
rect 222 -2672 278 -2580
rect 2350 -2672 2406 -2580
rect -3056 -3650 -3054 -2874
rect -3054 -3650 -3002 -2874
rect -3002 -3650 -3000 -2874
rect -2608 -3650 -2606 -2874
rect -2606 -3650 -2554 -2874
rect -2554 -3650 -2552 -2874
rect -2162 -3646 -2160 -2874
rect -2160 -3646 -2108 -2874
rect -2108 -3646 -2106 -2874
rect -1992 -3646 -1990 -2874
rect -1990 -3646 -1938 -2874
rect -1938 -3646 -1936 -2874
rect -1544 -3650 -1542 -2874
rect -1542 -3650 -1490 -2874
rect -1490 -3650 -1488 -2874
rect -1098 -3650 -1096 -2874
rect -1096 -3650 -1044 -2874
rect -1044 -3650 -1042 -2874
rect -928 -3648 -926 -2874
rect -926 -3648 -874 -2874
rect -874 -3648 -872 -2874
rect -480 -3650 -478 -2874
rect -478 -3650 -426 -2874
rect -426 -3650 -424 -2874
rect 222 -3136 276 -2948
rect 276 -3136 278 -2948
rect 986 -3136 988 -2948
rect 988 -3136 1040 -2948
rect 1040 -3136 1042 -2948
rect 2350 -3136 2404 -2948
rect 2404 -3136 2406 -2948
rect 3114 -3136 3116 -2948
rect 3116 -3136 3168 -2948
rect 3168 -3136 3170 -2948
rect 1812 -3556 1868 -3464
rect -3222 -4396 -3166 -4284
rect -1988 -4396 -1932 -4284
rect 1812 -4866 1814 -3890
rect 1814 -4866 1866 -3890
rect 1866 -4866 1868 -3890
<< metal3 >>
rect -2614 48 -2546 58
rect -2614 -394 -2608 48
rect -2552 -394 -2546 48
rect -3232 -1320 -3164 -1314
rect -3232 -2096 -3226 -1320
rect -3170 -2096 -3164 -1320
rect -3232 -2580 -3164 -2096
rect -3232 -2672 -3226 -2580
rect -3170 -2672 -3164 -2580
rect -3232 -4274 -3164 -2672
rect -3062 -1318 -2994 -1312
rect -3062 -2096 -3056 -1318
rect -3000 -2096 -2994 -1318
rect -3062 -2436 -2994 -2096
rect -3062 -2528 -3056 -2436
rect -3000 -2528 -2994 -2436
rect -3062 -2874 -2994 -2528
rect -3062 -3650 -3056 -2874
rect -3000 -3650 -2994 -2874
rect -3062 -3656 -2994 -3650
rect -2614 -1320 -2546 -394
rect -1550 48 -1482 58
rect -1550 -394 -1544 48
rect -1488 -394 -1482 48
rect -2614 -2096 -2608 -1320
rect -2552 -2096 -2546 -1320
rect -2614 -2874 -2546 -2096
rect -2614 -3650 -2608 -2874
rect -2552 -3650 -2546 -2874
rect -2614 -3656 -2546 -3650
rect -2168 -1318 -2100 -1312
rect -2168 -2090 -2162 -1318
rect -2106 -2090 -2100 -1318
rect -2168 -2436 -2100 -2090
rect -2168 -2528 -2162 -2436
rect -2106 -2528 -2100 -2436
rect -2168 -2874 -2100 -2528
rect -2168 -3646 -2162 -2874
rect -2106 -3646 -2100 -2874
rect -2168 -3652 -2100 -3646
rect -1998 -1318 -1930 -1312
rect -1998 -2096 -1992 -1318
rect -1936 -2096 -1930 -1318
rect -1998 -2436 -1930 -2096
rect -1998 -2528 -1992 -2436
rect -1936 -2528 -1930 -2436
rect -1998 -2874 -1930 -2528
rect -1998 -3646 -1992 -2874
rect -1936 -3646 -1930 -2874
rect -1998 -4274 -1930 -3646
rect -1550 -1320 -1482 -394
rect -486 48 -418 58
rect -486 -394 -480 48
rect -424 -394 -418 48
rect -1550 -2096 -1544 -1320
rect -1488 -2096 -1482 -1320
rect -1550 -2874 -1482 -2096
rect -1550 -3650 -1544 -2874
rect -1488 -3650 -1482 -2874
rect -1550 -3656 -1482 -3650
rect -1104 -1318 -1036 -1312
rect -1104 -2090 -1098 -1318
rect -1042 -2090 -1036 -1318
rect -1104 -2436 -1036 -2090
rect -1104 -2528 -1098 -2436
rect -1042 -2528 -1036 -2436
rect -1104 -2874 -1036 -2528
rect -1104 -3650 -1098 -2874
rect -1042 -3650 -1036 -2874
rect -1104 -3656 -1036 -3650
rect -934 -1318 -866 -1312
rect -934 -2096 -928 -1318
rect -872 -2096 -866 -1318
rect -934 -2436 -866 -2096
rect -934 -2528 -928 -2436
rect -872 -2528 -866 -2436
rect -934 -2874 -866 -2528
rect -934 -3648 -928 -2874
rect -872 -3648 -866 -2874
rect -934 -3654 -866 -3648
rect -486 -1320 -418 -394
rect -486 -2096 -480 -1320
rect -424 -2096 -418 -1320
rect -486 -2874 -418 -2096
rect -486 -3650 -480 -2874
rect -424 -3650 -418 -2874
rect 216 -1320 284 -1314
rect 216 -2296 222 -1320
rect 278 -2296 284 -1320
rect 216 -2580 284 -2296
rect 2344 -1320 2412 -1314
rect 2344 -2296 2350 -1320
rect 2406 -2296 2412 -1320
rect 978 -2344 1050 -2338
rect 978 -2400 984 -2344
rect 1044 -2400 1050 -2344
rect 978 -2406 1050 -2400
rect 216 -2672 222 -2580
rect 278 -2672 284 -2580
rect 216 -2948 284 -2672
rect 216 -3136 222 -2948
rect 278 -3136 284 -2948
rect 216 -3146 284 -3136
rect 980 -2948 1048 -2406
rect 980 -3136 986 -2948
rect 1042 -3136 1048 -2948
rect 980 -3146 1048 -3136
rect 2344 -2580 2412 -2296
rect 3106 -2342 3178 -2336
rect 3106 -2398 3112 -2342
rect 3172 -2398 3178 -2342
rect 3106 -2404 3178 -2398
rect 2344 -2672 2350 -2580
rect 2406 -2672 2412 -2580
rect 2344 -2948 2412 -2672
rect 2344 -3136 2350 -2948
rect 2406 -3136 2412 -2948
rect 2344 -3146 2412 -3136
rect 3108 -2948 3176 -2404
rect 3108 -3136 3114 -2948
rect 3170 -3136 3176 -2948
rect 3108 -3146 3176 -3136
rect -486 -3656 -418 -3650
rect 1806 -3464 1874 -3458
rect 1806 -3556 1812 -3464
rect 1868 -3556 1874 -3464
rect 1806 -3890 1874 -3556
rect -3232 -4284 -3160 -4274
rect -3232 -4396 -3222 -4284
rect -3166 -4396 -3160 -4284
rect -3232 -4406 -3160 -4396
rect -1998 -4284 -1926 -4274
rect -1998 -4396 -1988 -4284
rect -1932 -4396 -1926 -4284
rect -1998 -4406 -1926 -4396
rect 1806 -4866 1812 -3890
rect 1868 -4866 1874 -3890
rect 1806 -4872 1874 -4866
use sky130_fd_pr__pfet_01v8_lvt_AGRSB2  M4
timestamp 1682091667
transform 1 0 -4036 0 1 -1730
box -294 -264 294 298
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M5
timestamp 1681340463
transform -1 0 -3416 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__pfet_01v8_lvt_AGRSB2  M12
timestamp 1682091667
transform 1 0 -4946 0 -1 -1696
box -294 -264 294 298
use sky130_fd_pr__pfet_01v8_lvt_AGRSB2  M13
timestamp 1682091667
transform -1 0 -5552 0 -1 -1696
box -294 -264 294 298
use sky130_fd_pr__pfet_01v8_lvt_AGRSB2  M14
timestamp 1682091667
transform 1 0 -4946 0 -1 -2512
box -294 -264 294 298
use sky130_fd_pr__pfet_01v8_lvt_AGRSB2  M15
timestamp 1682091667
transform -1 0 -5552 0 -1 -2512
box -294 -264 294 298
use sky130_fd_pr__nfet_01v8_lvt_69Y42S  M16
timestamp 1682094193
transform 1 0 -4946 0 1 -2979
box -258 -107 258 107
use sky130_fd_pr__nfet_01v8_lvt_69Y42S  M17
timestamp 1682094193
transform -1 0 -5552 0 1 -2979
box -258 -107 258 107
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M61
timestamp 1681340463
transform 1 0 -2810 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M62
timestamp 1681340463
transform 1 0 -2352 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M63
timestamp 1681340463
transform -1 0 -1746 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M64
timestamp 1681340463
transform 1 0 -1288 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_P3X5Q9  M65
timestamp 1681340463
transform 1 0 -682 0 1 -1739
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M66
timestamp 1681340463
transform 1 0 -2810 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M67
timestamp 1681340463
transform 1 0 -2352 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M68
timestamp 1681340463
transform 1 0 -1746 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M69
timestamp 1681340463
transform 1 0 -1288 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__nfet_01v8_lvt_N4YUK3  M71
timestamp 1682091667
transform 1 0 786 0 1 -3005
box -258 -157 258 157
use sky130_fd_pr__nfet_01v8_lvt_N4YUK3  M72
timestamp 1682091667
transform 1 0 1244 0 1 -3005
box -258 -157 258 157
use sky130_fd_pr__nfet_01v8_lvt_N4YUK3  M73
timestamp 1682091667
transform 1 0 2914 0 1 -3005
box -258 -157 258 157
use sky130_fd_pr__nfet_01v8_lvt_N4YUK3  M74
timestamp 1682091667
transform 1 0 3372 0 1 -3005
box -258 -157 258 157
use sky130_fd_pr__nfet_01v8_lvt_ULR8M5  M81
timestamp 1682091667
transform 1 0 172 0 1 -3005
box -108 -157 108 157
use sky130_fd_pr__nfet_01v8_lvt_ULR8M5  M82
timestamp 1682091667
transform 1 0 330 0 1 -3005
box -108 -157 108 157
use sky130_fd_pr__nfet_01v8_lvt_ULR8M5  M83
timestamp 1682091667
transform 1 0 2300 0 1 -3005
box -108 -157 108 157
use sky130_fd_pr__nfet_01v8_lvt_ULR8M5  M84
timestamp 1682091667
transform 1 0 2458 0 1 -3005
box -108 -157 108 157
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M91
timestamp 1681382244
transform 1 0 3214 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M92
timestamp 1681382244
transform 1 0 3672 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M93
timestamp 1681382244
transform 1 0 1086 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M94
timestamp 1681382244
transform 1 0 1544 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M101
timestamp 1681382244
transform 1 0 22 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M102
timestamp 1681382244
transform 1 0 480 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M103
timestamp 1681382244
transform 1 0 2150 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__pfet_01v8_lvt_HLJ7ZV  M104
timestamp 1681382244
transform 1 0 2608 0 1 -1844
box -294 -564 294 598
use sky130_fd_pr__nfet_01v8_D8YEEC  M111
timestamp 1681382244
transform 1 0 1006 0 1 -4349
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_D8YEEC  M112
timestamp 1681382244
transform 1 0 1612 0 1 -4349
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_D8YEEC  M113
timestamp 1681382244
transform 1 0 2070 0 1 -4349
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_D8YEEC  M114
timestamp 1681382244
transform 1 0 2676 0 1 -4349
box -258 -557 258 557
use sky130_fd_pr__nfet_01v8_lvt_69YEWK  M610
timestamp 1681340463
transform 1 0 -682 0 1 -3231
box -258 -457 258 457
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q3 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1671334046
transform 1 0 -3018 0 1 -4738
box 0 0 796 796
use sky130_fd_pr__pnp_05v5_W3p40L3p40  Q4
timestamp 1671334046
transform 1 0 -1824 0 1 -4738
box 0 0 796 796
<< labels >>
flabel metal2 -5848 -5776 4348 -5308 0 FreeMono 1920 0 0 0 vss
port 0 nsew
flabel metal2 -5848 -404 4348 64 0 FreeMono 1920 0 0 0 vdd
port 1 nsew
flabel metal1 4174 -4880 4348 -4080 0 FreeMono 960 90 0 0 vtemp
port 2 nsew
<< end >>
