* NGSPICE file created from Temperature_Sensor.ext - technology: sky130A

.subckt Temperature_Sensor vtemp vdd vss
M610 a_n3070_n3662# a_n3836_n1894# vdd vss sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=8.6 as=0.58 ps=4.29 w=4 l=2
M69 a_n3070_n3662# a_n3836_n1894# vdd vss sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=8.6 as=0.58 ps=4.29 w=4 l=2
M15 a_n5752_n3086# a_n5752_n2774# a_n5810_n2748# vdd sky130_fd_pr__pfet_01v8_lvt ad=0.6 pd=4.6 as=0.58 ps=4.58 w=2 l=2
M91 a_n178_n2405# a_n178_n2405# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=1.5 ps=10.6 w=5 l=2
M5 a_n3216_n2108# a_n3836_n1894# a_n3836_n1894# vss sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=8.6 as=1.16 ps=8.58 w=4 l=2
M92 vdd a_n178_n2405# a_n178_n2405# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.6 as=0.725 ps=5.29 w=5 l=2
M68 vdd a_n3836_n1894# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.2 ps=8.6 w=4 l=2
M93 a_n178_n2405# a_n178_n2405# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=1.5 ps=10.6 w=5 l=2
M16 vss a_n5752_n2774# a_n5752_n2774# vss sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.58 as=0.15 ps=1.6 w=0.5 l=2
M81 vtemp a_n3070_n3662# a_62_n3136# vss sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.3 ps=2.6 w=1 l=0.5
M71 a_62_n3136# a_n3216_n2108# a_n178_n2405# vss sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.145 ps=1.29 w=1 l=2
M67 vdd a_n3836_n1894# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.2 ps=8.6 w=4 l=2
M111 vss a_n5752_n2774# a_62_n3136# vss sky130_fd_pr__nfet_01v8 ad=1.5 pd=10.6 as=1.45 ps=10.6 w=5 l=2
M112 vss a_n5752_n2774# a_62_n3136# vss sky130_fd_pr__nfet_01v8 ad=1.5 pd=10.6 as=0.725 ps=5.29 w=5 l=2
Q3 vss vss a_n3216_n2108# sky130_fd_pr__pnp_05v5_W3p40L3p40
M12 a_n5752_n1958# a_n5752_n1958# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.6 ps=4.6 w=2 l=2
M66 vdd a_n3836_n1894# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.2 ps=8.6 w=4 l=2
M65 a_n3070_n3662# a_n3836_n1894# vdd vss sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=8.6 as=0.58 ps=4.29 w=4 l=2
Q4 vss vss a_n3070_n3662# sky130_fd_pr__pnp_05v5_W3p40L3p40
M72 a_62_n3136# a_n3216_n2108# a_n178_n2405# vss sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.145 ps=1.29 w=1 l=2
M113 a_62_n3136# a_n5752_n2774# vss vss sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.5 ps=10.6 w=5 l=2
M101 vdd a_n178_n2405# vtemp vdd sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.6 as=0.725 ps=5.29 w=5 l=2
M102 vtemp a_n178_n2405# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=1.5 ps=10.6 w=5 l=2
M82 vtemp a_n3070_n3662# a_62_n3136# vss sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.3 ps=2.6 w=1 l=0.5
M73 a_n178_n2405# a_n3216_n2108# a_62_n3136# vss sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.3 ps=2.6 w=1 l=2
M74 a_n178_n2405# a_n3216_n2108# a_62_n3136# vss sky130_fd_pr__nfet_01v8_lvt ad=0.145 pd=1.29 as=0.3 ps=2.6 w=1 l=2
M64 a_n3070_n3662# a_n3836_n1894# vdd vss sky130_fd_pr__nfet_01v8_lvt ad=1.2 pd=8.6 as=0.58 ps=4.29 w=4 l=2
M4 a_n3836_n1894# a_n5752_n2774# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.6 ps=4.6 w=2 l=2
M14 a_n5752_n1958# a_n5752_n2774# a_n5752_n2774# vdd sky130_fd_pr__pfet_01v8_lvt ad=0.58 pd=4.58 as=0.6 ps=4.6 w=2 l=2
M17 a_n5752_n3086# a_n5752_n3086# vss vss sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.145 ps=1.58 w=0.5 l=2
M83 a_62_n3136# a_n3070_n3662# vtemp vss sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.145 ps=1.29 w=1 l=0.5
M63 vdd a_n3836_n1894# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.2 ps=8.6 w=4 l=2
M62 vdd a_n3836_n1894# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=0.58 pd=4.29 as=1.2 ps=8.6 w=4 l=2
M13 vdd a_n5752_n1958# a_n5810_n2748# vdd sky130_fd_pr__pfet_01v8_lvt ad=0.6 pd=4.6 as=0.58 ps=4.58 w=2 l=2
M103 vtemp a_n178_n2405# vdd vdd sky130_fd_pr__pfet_01v8_lvt ad=0.725 pd=5.29 as=1.5 ps=10.6 w=5 l=2
M114 a_62_n3136# a_n5752_n2774# vss vss sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.5 ps=10.6 w=5 l=2
M104 vdd a_n178_n2405# vtemp vdd sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.6 as=0.725 ps=5.29 w=5 l=2
M94 vdd a_n178_n2405# a_n178_n2405# vdd sky130_fd_pr__pfet_01v8_lvt ad=1.5 pd=10.6 as=0.725 ps=5.29 w=5 l=2
M84 a_62_n3136# a_n3070_n3662# vtemp vss sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.6 as=0.145 ps=1.29 w=1 l=0.5
M61 vdd a_n3836_n1894# a_n3070_n3662# vss sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.2 ps=8.6 w=4 l=2
.ends

