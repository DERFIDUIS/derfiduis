** sch_path: /home/karlajcm/Documentos/TESIS DE
*+ GRADO/WORK_IN_PROGRESS/My_xschem/ring_oscillator_tb.sch
**.subckt ring_oscillator_tb vosc vdd vtemp
*.iopin vosc
*.iopin vdd
*.iopin vtemp
Vdd vdd GND 1.5
.save i(vdd)
vtemp vtemp GND 0.01
.save i(vtemp)
x1 vtemp vosc GND vdd ring_oscillator
**** begin user architecture code

.control
save all
nodeset v(vosc)=0


let v_xmax= 1.81
let step= 0.01
let v_x = 0
let i=0


* These vector will be used to save the data of each iteration.
let freqs = unitvec(180)
let volts = unitvec(180)

* Start loop
while v_x <= v_xmax

* Modify Vtemp
  alter vtemp = v_x

* Run transient analysis
  tran 2.5n 500n 

* Find period 
  echo
  meas  TRAN  period  TRIG  v(vosc) VAL=1.2 RISE=20  TARG v(vosc)  VAL=1.2 RISE=21
  echo


* Save freq and vtemp in vectors
  let freqs[i] = 1/period
  let volts[i] = v_x

* Modify widths
  let v_x = v_x + step
  
 * Counter increment
  let i = i + 1
  	
end
  plot vosc
* Export vector data into raw file
write ring_oscilator_tb.raw freqs volts

* Plot frequency vs Vtemp
  plot freqs vs volts

.endc


** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /usr/local/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

.include ring_oscillator.spice

.GLOBAL GND
.end
