** sch_path: /home/karlajcm/Documentos/TESIS DE
*+ GRADO/WORK_IN_PROGRESS/My_xschem/For_Layout/OPAMP_lvt_PMOS.sch
.subckt OPAMP_lvt_PMOS vdd vss out vinp vinn
*.PININFO vdd:B vss:B out:B vinp:B vinn:B
XC2 net3 out sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
M11 net1 net4 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M21 net2 vinn net1 vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M31 net3 vinp net1 vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M41 net2 net2 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
M51 net3 net2 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
M61 out net4 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M71 out net3 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
M81 net4 net4 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M91 net4 net4 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
M92 net4 net4 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
M82 net4 net4 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M12 net1 net4 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M22 net2 vinn net1 vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M23 net2 vinn net1 vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M24 net2 vinn net1 vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M42 net2 net2 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
M34 net3 vinp net1 vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M33 net3 vinp net1 vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M32 net3 vinp net1 vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M52 net3 net2 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
M62 out net4 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=5 nf=1 m=1
M72 out net3 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
M73 out net3 vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=2 nf=1 m=1
.ends
.end
