magic
tech sky130A
timestamp 1682034855
<< metal4 >>
rect -448337 52271 -444394 52283
rect -447983 43844 -444394 52271
rect -441548 52271 -437605 52283
rect -441548 43844 -437959 52271
rect -447983 35777 -444240 43844
rect -441591 35777 -437959 43844
rect -447983 27295 -444394 35777
rect -448337 27283 -444394 27295
rect -441548 27295 -437959 35777
rect -441548 27283 -437605 27295
<< via4 >>
rect -448337 27295 -447983 52271
rect -437959 27295 -437605 52271
<< metal5 >>
rect -586971 350283 -298971 375283
rect -586971 52283 -561971 350283
rect -323971 52283 -298971 350283
rect -586971 52271 -447971 52283
rect -586971 27295 -448337 52271
rect -447983 27295 -447971 52271
rect -586971 27283 -447971 27295
rect -437971 52271 -298971 52283
rect -437971 27295 -437959 52271
rect -437605 27295 -298971 52271
rect -437971 27283 -298971 27295
use sky130_fd_pr__cap_mim_m3_1_JMY65W  sky130_fd_pr__cap_mim_m3_1_JMY65W_0
timestamp 1682034855
transform 1 0 -442935 0 1 42531
box -1373 -1300 1373 1300
use sky130_fd_pr__cap_mim_m3_1_JMY65W  sky130_fd_pr__cap_mim_m3_1_JMY65W_1
timestamp 1682034855
transform 1 0 -442929 0 1 39811
box -1373 -1300 1373 1300
use sky130_fd_pr__cap_mim_m3_1_UXZFBW  sky130_fd_pr__cap_mim_m3_1_UXZFBW_0
timestamp 1682034855
transform 1 0 -442928 0 1 37090
box -1373 -1301 1373 1301
<< end >>
