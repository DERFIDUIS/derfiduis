magic
tech sky130A
magscale 1 2
timestamp 1681576725
<< error_p >>
rect -758 -531 -700 469
rect 700 -531 758 469
<< nmoslvt >>
rect -700 -531 700 469
<< ndiff >>
rect -758 457 -700 469
rect -758 -519 -746 457
rect -712 -519 -700 457
rect -758 -531 -700 -519
rect 700 457 758 469
rect 700 -519 712 457
rect 746 -519 758 457
rect 700 -531 758 -519
<< ndiffc >>
rect -746 -519 -712 457
rect 712 -519 746 457
<< poly >>
rect -700 541 700 557
rect -700 507 -684 541
rect 684 507 700 541
rect -700 469 700 507
rect -700 -557 700 -531
<< polycont >>
rect -684 507 684 541
<< locali >>
rect -700 507 -684 541
rect 684 507 700 541
rect -746 457 -712 473
rect -746 -535 -712 -519
rect 712 457 746 473
rect 712 -535 746 -519
<< viali >>
rect -684 507 684 541
rect -746 -519 -712 457
rect 712 -519 746 457
<< metal1 >>
rect -696 541 696 547
rect -696 507 -684 541
rect 684 507 696 541
rect -696 501 696 507
rect -752 457 -706 469
rect -752 -519 -746 457
rect -712 -519 -706 457
rect -752 -531 -706 -519
rect 706 457 752 469
rect 706 -519 712 457
rect 746 -519 752 457
rect 706 -531 752 -519
<< properties >>
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.0 l 7.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
