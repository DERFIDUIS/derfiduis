magic
tech sky130A
magscale 1 2
timestamp 1681769244
<< nwell >>
rect 3458 -2414 3572 -652
rect 4534 -2414 4636 -652
rect 2852 -2868 2918 -2748
rect 2852 -2902 2926 -2868
rect 2852 -2936 2918 -2902
rect 2852 -2970 2926 -2936
rect 2852 -3004 2918 -2970
rect 2852 -3038 2926 -3004
rect 2852 -3072 2918 -3038
rect 2852 -3106 2926 -3072
rect 2852 -3140 2918 -3106
rect 2852 -3174 2926 -3140
rect 2852 -3208 2918 -3174
rect 2852 -3242 2926 -3208
rect 2852 -3276 2918 -3242
rect 2852 -3310 2926 -3276
rect 2852 -3344 2918 -3310
rect 2852 -3378 2926 -3344
rect 2852 -3412 2918 -3378
rect 2852 -3446 2926 -3412
rect 2852 -3480 2918 -3446
rect 2852 -3514 2926 -3480
rect 2852 -3710 2918 -3514
rect 3990 -3710 4104 -2748
<< pwell >>
rect 546 -7834 782 -4150
rect 1152 -7834 1388 -4150
rect 1758 -7832 1994 -4148
rect 2004 -4572 2252 -4570
rect 2364 -7832 2600 -4148
rect 2970 -7832 3206 -4148
rect 3576 -7832 3812 -4148
rect 4182 -7832 4418 -4148
rect 4788 -7832 5024 -4148
rect 5394 -7832 5630 -4148
rect 6000 -7832 6236 -4148
<< pdiff >>
rect 3470 -2314 3472 -714
rect 3558 -2314 3560 -714
rect 4534 -2314 4536 -714
rect 2952 -3610 2954 -2810
rect 4002 -3610 4004 -2810
rect 4090 -3610 4092 -2810
<< psubdiff >>
rect 546 -4166 674 -4150
rect 546 -4338 570 -4166
rect 650 -4338 674 -4166
rect 546 -4510 674 -4338
rect 546 -4682 570 -4510
rect 650 -4682 674 -4510
rect 546 -4854 674 -4682
rect 546 -5026 570 -4854
rect 650 -5026 674 -4854
rect 546 -5198 674 -5026
rect 546 -5370 570 -5198
rect 650 -5370 674 -5198
rect 546 -5542 674 -5370
rect 546 -5714 570 -5542
rect 650 -5714 674 -5542
rect 546 -5886 674 -5714
rect 546 -6058 570 -5886
rect 650 -6058 674 -5886
rect 546 -6230 674 -6058
rect 546 -6402 570 -6230
rect 650 -6402 674 -6230
rect 546 -6574 674 -6402
rect 546 -6746 570 -6574
rect 650 -6746 674 -6574
rect 546 -6918 674 -6746
rect 546 -7090 570 -6918
rect 650 -7090 674 -6918
rect 546 -7262 674 -7090
rect 546 -7434 570 -7262
rect 650 -7434 674 -7262
rect 546 -7606 674 -7434
rect 546 -7778 570 -7606
rect 650 -7778 674 -7606
rect 546 -7834 674 -7778
rect 1152 -4166 1280 -4150
rect 1152 -4338 1176 -4166
rect 1256 -4338 1280 -4166
rect 1152 -4510 1280 -4338
rect 1152 -4682 1176 -4510
rect 1256 -4682 1280 -4510
rect 1152 -4854 1280 -4682
rect 1152 -5026 1176 -4854
rect 1256 -5026 1280 -4854
rect 1152 -5198 1280 -5026
rect 1152 -5370 1176 -5198
rect 1256 -5370 1280 -5198
rect 1152 -5542 1280 -5370
rect 1152 -5714 1176 -5542
rect 1256 -5714 1280 -5542
rect 1152 -5886 1280 -5714
rect 1152 -6058 1176 -5886
rect 1256 -6058 1280 -5886
rect 1152 -6230 1280 -6058
rect 1152 -6402 1176 -6230
rect 1256 -6402 1280 -6230
rect 1152 -6574 1280 -6402
rect 1152 -6746 1176 -6574
rect 1256 -6746 1280 -6574
rect 1152 -6918 1280 -6746
rect 1152 -7090 1176 -6918
rect 1256 -7090 1280 -6918
rect 1152 -7262 1280 -7090
rect 1152 -7434 1176 -7262
rect 1256 -7434 1280 -7262
rect 1152 -7606 1280 -7434
rect 1152 -7778 1176 -7606
rect 1256 -7778 1280 -7606
rect 1152 -7834 1280 -7778
rect 1758 -4164 1886 -4148
rect 1758 -4336 1782 -4164
rect 1862 -4336 1886 -4164
rect 1758 -4508 1886 -4336
rect 1758 -4680 1782 -4508
rect 1862 -4680 1886 -4508
rect 1758 -4852 1886 -4680
rect 1758 -5024 1782 -4852
rect 1862 -5024 1886 -4852
rect 1758 -5196 1886 -5024
rect 1758 -5368 1782 -5196
rect 1862 -5368 1886 -5196
rect 1758 -5540 1886 -5368
rect 1758 -5712 1782 -5540
rect 1862 -5712 1886 -5540
rect 1758 -5884 1886 -5712
rect 1758 -6056 1782 -5884
rect 1862 -6056 1886 -5884
rect 1758 -6228 1886 -6056
rect 1758 -6400 1782 -6228
rect 1862 -6400 1886 -6228
rect 1758 -6572 1886 -6400
rect 1758 -6744 1782 -6572
rect 1862 -6744 1886 -6572
rect 1758 -6916 1886 -6744
rect 1758 -7088 1782 -6916
rect 1862 -7088 1886 -6916
rect 1758 -7260 1886 -7088
rect 1758 -7432 1782 -7260
rect 1862 -7432 1886 -7260
rect 1758 -7604 1886 -7432
rect 1758 -7776 1782 -7604
rect 1862 -7776 1886 -7604
rect 1758 -7832 1886 -7776
rect 2364 -4164 2492 -4148
rect 2364 -4336 2388 -4164
rect 2468 -4336 2492 -4164
rect 2364 -4508 2492 -4336
rect 2364 -4680 2388 -4508
rect 2468 -4680 2492 -4508
rect 2364 -4852 2492 -4680
rect 2364 -5024 2388 -4852
rect 2468 -5024 2492 -4852
rect 2364 -5196 2492 -5024
rect 2364 -5368 2388 -5196
rect 2468 -5368 2492 -5196
rect 2364 -5540 2492 -5368
rect 2364 -5712 2388 -5540
rect 2468 -5712 2492 -5540
rect 2364 -5884 2492 -5712
rect 2364 -6056 2388 -5884
rect 2468 -6056 2492 -5884
rect 2364 -6228 2492 -6056
rect 2364 -6400 2388 -6228
rect 2468 -6400 2492 -6228
rect 2364 -6572 2492 -6400
rect 2364 -6744 2388 -6572
rect 2468 -6744 2492 -6572
rect 2364 -6916 2492 -6744
rect 2364 -7088 2388 -6916
rect 2468 -7088 2492 -6916
rect 2364 -7260 2492 -7088
rect 2364 -7432 2388 -7260
rect 2468 -7432 2492 -7260
rect 2364 -7604 2492 -7432
rect 2364 -7776 2388 -7604
rect 2468 -7776 2492 -7604
rect 2364 -7832 2492 -7776
rect 2970 -4164 3098 -4148
rect 2970 -4336 2994 -4164
rect 3074 -4336 3098 -4164
rect 2970 -4508 3098 -4336
rect 2970 -4680 2994 -4508
rect 3074 -4680 3098 -4508
rect 2970 -4852 3098 -4680
rect 2970 -5024 2994 -4852
rect 3074 -5024 3098 -4852
rect 2970 -5196 3098 -5024
rect 2970 -5368 2994 -5196
rect 3074 -5368 3098 -5196
rect 2970 -5540 3098 -5368
rect 2970 -5712 2994 -5540
rect 3074 -5712 3098 -5540
rect 2970 -5884 3098 -5712
rect 2970 -6056 2994 -5884
rect 3074 -6056 3098 -5884
rect 2970 -6228 3098 -6056
rect 2970 -6400 2994 -6228
rect 3074 -6400 3098 -6228
rect 2970 -6572 3098 -6400
rect 2970 -6744 2994 -6572
rect 3074 -6744 3098 -6572
rect 2970 -6916 3098 -6744
rect 2970 -7088 2994 -6916
rect 3074 -7088 3098 -6916
rect 2970 -7260 3098 -7088
rect 2970 -7432 2994 -7260
rect 3074 -7432 3098 -7260
rect 2970 -7604 3098 -7432
rect 2970 -7776 2994 -7604
rect 3074 -7776 3098 -7604
rect 2970 -7832 3098 -7776
rect 3576 -4164 3704 -4148
rect 3576 -4336 3600 -4164
rect 3680 -4336 3704 -4164
rect 3576 -4508 3704 -4336
rect 3576 -4680 3600 -4508
rect 3680 -4680 3704 -4508
rect 3576 -4852 3704 -4680
rect 3576 -5024 3600 -4852
rect 3680 -5024 3704 -4852
rect 3576 -5196 3704 -5024
rect 3576 -5368 3600 -5196
rect 3680 -5368 3704 -5196
rect 3576 -5540 3704 -5368
rect 3576 -5712 3600 -5540
rect 3680 -5712 3704 -5540
rect 3576 -5884 3704 -5712
rect 3576 -6056 3600 -5884
rect 3680 -6056 3704 -5884
rect 3576 -6228 3704 -6056
rect 3576 -6400 3600 -6228
rect 3680 -6400 3704 -6228
rect 3576 -6572 3704 -6400
rect 3576 -6744 3600 -6572
rect 3680 -6744 3704 -6572
rect 3576 -6916 3704 -6744
rect 3576 -7088 3600 -6916
rect 3680 -7088 3704 -6916
rect 3576 -7260 3704 -7088
rect 3576 -7432 3600 -7260
rect 3680 -7432 3704 -7260
rect 3576 -7604 3704 -7432
rect 3576 -7776 3600 -7604
rect 3680 -7776 3704 -7604
rect 3576 -7832 3704 -7776
rect 4182 -4164 4310 -4148
rect 4182 -4336 4206 -4164
rect 4286 -4336 4310 -4164
rect 4182 -4508 4310 -4336
rect 4182 -4680 4206 -4508
rect 4286 -4680 4310 -4508
rect 4182 -4852 4310 -4680
rect 4182 -5024 4206 -4852
rect 4286 -5024 4310 -4852
rect 4182 -5196 4310 -5024
rect 4182 -5368 4206 -5196
rect 4286 -5368 4310 -5196
rect 4182 -5540 4310 -5368
rect 4182 -5712 4206 -5540
rect 4286 -5712 4310 -5540
rect 4182 -5884 4310 -5712
rect 4182 -6056 4206 -5884
rect 4286 -6056 4310 -5884
rect 4182 -6228 4310 -6056
rect 4182 -6400 4206 -6228
rect 4286 -6400 4310 -6228
rect 4182 -6572 4310 -6400
rect 4182 -6744 4206 -6572
rect 4286 -6744 4310 -6572
rect 4182 -6916 4310 -6744
rect 4182 -7088 4206 -6916
rect 4286 -7088 4310 -6916
rect 4182 -7260 4310 -7088
rect 4182 -7432 4206 -7260
rect 4286 -7432 4310 -7260
rect 4182 -7604 4310 -7432
rect 4182 -7776 4206 -7604
rect 4286 -7776 4310 -7604
rect 4182 -7832 4310 -7776
rect 4788 -4164 4916 -4148
rect 4788 -4336 4812 -4164
rect 4892 -4336 4916 -4164
rect 4788 -4508 4916 -4336
rect 4788 -4680 4812 -4508
rect 4892 -4680 4916 -4508
rect 4788 -4852 4916 -4680
rect 4788 -5024 4812 -4852
rect 4892 -5024 4916 -4852
rect 4788 -5196 4916 -5024
rect 4788 -5368 4812 -5196
rect 4892 -5368 4916 -5196
rect 4788 -5540 4916 -5368
rect 4788 -5712 4812 -5540
rect 4892 -5712 4916 -5540
rect 4788 -5884 4916 -5712
rect 4788 -6056 4812 -5884
rect 4892 -6056 4916 -5884
rect 4788 -6228 4916 -6056
rect 4788 -6400 4812 -6228
rect 4892 -6400 4916 -6228
rect 4788 -6572 4916 -6400
rect 4788 -6744 4812 -6572
rect 4892 -6744 4916 -6572
rect 4788 -6916 4916 -6744
rect 4788 -7088 4812 -6916
rect 4892 -7088 4916 -6916
rect 4788 -7260 4916 -7088
rect 4788 -7432 4812 -7260
rect 4892 -7432 4916 -7260
rect 4788 -7604 4916 -7432
rect 4788 -7776 4812 -7604
rect 4892 -7776 4916 -7604
rect 4788 -7832 4916 -7776
rect 5394 -4164 5522 -4148
rect 5394 -4336 5418 -4164
rect 5498 -4336 5522 -4164
rect 5394 -4508 5522 -4336
rect 5394 -4680 5418 -4508
rect 5498 -4680 5522 -4508
rect 5394 -4852 5522 -4680
rect 5394 -5024 5418 -4852
rect 5498 -5024 5522 -4852
rect 5394 -5196 5522 -5024
rect 5394 -5368 5418 -5196
rect 5498 -5368 5522 -5196
rect 5394 -5540 5522 -5368
rect 5394 -5712 5418 -5540
rect 5498 -5712 5522 -5540
rect 5394 -5884 5522 -5712
rect 5394 -6056 5418 -5884
rect 5498 -6056 5522 -5884
rect 5394 -6228 5522 -6056
rect 5394 -6400 5418 -6228
rect 5498 -6400 5522 -6228
rect 5394 -6572 5522 -6400
rect 5394 -6744 5418 -6572
rect 5498 -6744 5522 -6572
rect 5394 -6916 5522 -6744
rect 5394 -7088 5418 -6916
rect 5498 -7088 5522 -6916
rect 5394 -7260 5522 -7088
rect 5394 -7432 5418 -7260
rect 5498 -7432 5522 -7260
rect 5394 -7604 5522 -7432
rect 5394 -7776 5418 -7604
rect 5498 -7776 5522 -7604
rect 5394 -7832 5522 -7776
rect 6000 -4164 6128 -4148
rect 6000 -4336 6024 -4164
rect 6104 -4336 6128 -4164
rect 6000 -4508 6128 -4336
rect 6000 -4680 6024 -4508
rect 6104 -4680 6128 -4508
rect 6000 -4852 6128 -4680
rect 6000 -5024 6024 -4852
rect 6104 -5024 6128 -4852
rect 6000 -5196 6128 -5024
rect 6000 -5368 6024 -5196
rect 6104 -5368 6128 -5196
rect 6000 -5540 6128 -5368
rect 6000 -5712 6024 -5540
rect 6104 -5712 6128 -5540
rect 6000 -5884 6128 -5712
rect 6000 -6056 6024 -5884
rect 6104 -6056 6128 -5884
rect 6000 -6228 6128 -6056
rect 6000 -6400 6024 -6228
rect 6104 -6400 6128 -6228
rect 6000 -6572 6128 -6400
rect 6000 -6744 6024 -6572
rect 6104 -6744 6128 -6572
rect 6000 -6916 6128 -6744
rect 6000 -7088 6024 -6916
rect 6104 -7088 6128 -6916
rect 6000 -7260 6128 -7088
rect 6000 -7432 6024 -7260
rect 6104 -7432 6128 -7260
rect 6000 -7604 6128 -7432
rect 6000 -7776 6024 -7604
rect 6104 -7776 6128 -7604
rect 6000 -7832 6128 -7776
<< nsubdiff >>
rect 3472 -756 3558 -714
rect 3472 -790 3498 -756
rect 3532 -790 3558 -756
rect 3472 -824 3558 -790
rect 3472 -858 3498 -824
rect 3532 -858 3558 -824
rect 3472 -892 3558 -858
rect 3472 -926 3498 -892
rect 3532 -926 3558 -892
rect 3472 -960 3558 -926
rect 3472 -994 3498 -960
rect 3532 -994 3558 -960
rect 3472 -1028 3558 -994
rect 3472 -1062 3498 -1028
rect 3532 -1062 3558 -1028
rect 3472 -1096 3558 -1062
rect 3472 -1130 3498 -1096
rect 3532 -1130 3558 -1096
rect 3472 -1164 3558 -1130
rect 3472 -1198 3498 -1164
rect 3532 -1198 3558 -1164
rect 3472 -1232 3558 -1198
rect 3472 -1266 3498 -1232
rect 3532 -1266 3558 -1232
rect 3472 -1300 3558 -1266
rect 3472 -1334 3498 -1300
rect 3532 -1334 3558 -1300
rect 3472 -1368 3558 -1334
rect 3472 -1402 3498 -1368
rect 3532 -1402 3558 -1368
rect 3472 -1436 3558 -1402
rect 3472 -1470 3498 -1436
rect 3532 -1470 3558 -1436
rect 3472 -1504 3558 -1470
rect 3472 -1538 3498 -1504
rect 3532 -1538 3558 -1504
rect 3472 -1572 3558 -1538
rect 3472 -1606 3498 -1572
rect 3532 -1606 3558 -1572
rect 3472 -1640 3558 -1606
rect 3472 -1674 3498 -1640
rect 3532 -1674 3558 -1640
rect 3472 -1708 3558 -1674
rect 3472 -1742 3498 -1708
rect 3532 -1742 3558 -1708
rect 3472 -1776 3558 -1742
rect 3472 -1810 3498 -1776
rect 3532 -1810 3558 -1776
rect 3472 -1844 3558 -1810
rect 3472 -1878 3498 -1844
rect 3532 -1878 3558 -1844
rect 3472 -1912 3558 -1878
rect 3472 -1946 3498 -1912
rect 3532 -1946 3558 -1912
rect 3472 -1980 3558 -1946
rect 3472 -2014 3498 -1980
rect 3532 -2014 3558 -1980
rect 3472 -2048 3558 -2014
rect 3472 -2082 3498 -2048
rect 3532 -2082 3558 -2048
rect 3472 -2116 3558 -2082
rect 3472 -2150 3498 -2116
rect 3532 -2150 3558 -2116
rect 3472 -2184 3558 -2150
rect 3472 -2218 3498 -2184
rect 3532 -2218 3558 -2184
rect 3472 -2252 3558 -2218
rect 3472 -2286 3498 -2252
rect 3532 -2286 3558 -2252
rect 3472 -2314 3558 -2286
rect 4536 -756 4600 -714
rect 4536 -790 4562 -756
rect 4596 -790 4600 -756
rect 4536 -824 4600 -790
rect 4536 -858 4562 -824
rect 4596 -858 4600 -824
rect 4536 -892 4600 -858
rect 4536 -926 4562 -892
rect 4596 -926 4600 -892
rect 4536 -960 4600 -926
rect 4536 -994 4562 -960
rect 4596 -994 4600 -960
rect 4536 -1028 4600 -994
rect 4536 -1062 4562 -1028
rect 4596 -1062 4600 -1028
rect 4536 -1096 4600 -1062
rect 4536 -1130 4562 -1096
rect 4596 -1130 4600 -1096
rect 4536 -1164 4600 -1130
rect 4536 -1198 4562 -1164
rect 4596 -1198 4600 -1164
rect 4536 -1232 4600 -1198
rect 4536 -1266 4562 -1232
rect 4596 -1266 4600 -1232
rect 4536 -1300 4600 -1266
rect 4536 -1334 4562 -1300
rect 4596 -1334 4600 -1300
rect 4536 -1368 4600 -1334
rect 4536 -1402 4562 -1368
rect 4596 -1402 4600 -1368
rect 4536 -1436 4600 -1402
rect 4536 -1470 4562 -1436
rect 4596 -1470 4600 -1436
rect 4536 -1504 4600 -1470
rect 4536 -1538 4562 -1504
rect 4596 -1538 4600 -1504
rect 4536 -1572 4600 -1538
rect 4536 -1606 4562 -1572
rect 4596 -1606 4600 -1572
rect 4536 -1640 4600 -1606
rect 4536 -1674 4562 -1640
rect 4596 -1674 4600 -1640
rect 4536 -1708 4600 -1674
rect 4536 -1742 4562 -1708
rect 4596 -1742 4600 -1708
rect 4536 -1776 4600 -1742
rect 4536 -1810 4562 -1776
rect 4596 -1810 4600 -1776
rect 4536 -1844 4600 -1810
rect 4536 -1878 4562 -1844
rect 4596 -1878 4600 -1844
rect 4536 -1912 4600 -1878
rect 4536 -1946 4562 -1912
rect 4596 -1946 4600 -1912
rect 4536 -1980 4600 -1946
rect 4536 -2014 4562 -1980
rect 4596 -2014 4600 -1980
rect 4536 -2048 4600 -2014
rect 4536 -2082 4562 -2048
rect 4596 -2082 4600 -2048
rect 4536 -2116 4600 -2082
rect 4536 -2150 4562 -2116
rect 4596 -2150 4600 -2116
rect 4536 -2184 4600 -2150
rect 4536 -2218 4562 -2184
rect 4596 -2218 4600 -2184
rect 4536 -2252 4600 -2218
rect 4536 -2286 4562 -2252
rect 4596 -2286 4600 -2252
rect 4536 -2314 4600 -2286
rect 2888 -2868 2952 -2810
rect 2888 -2902 2892 -2868
rect 2926 -2902 2952 -2868
rect 2888 -2936 2952 -2902
rect 2888 -2970 2892 -2936
rect 2926 -2970 2952 -2936
rect 2888 -3004 2952 -2970
rect 2888 -3038 2892 -3004
rect 2926 -3038 2952 -3004
rect 2888 -3072 2952 -3038
rect 2888 -3106 2892 -3072
rect 2926 -3106 2952 -3072
rect 2888 -3140 2952 -3106
rect 2888 -3174 2892 -3140
rect 2926 -3174 2952 -3140
rect 2888 -3208 2952 -3174
rect 2888 -3242 2892 -3208
rect 2926 -3242 2952 -3208
rect 2888 -3276 2952 -3242
rect 2888 -3310 2892 -3276
rect 2926 -3310 2952 -3276
rect 2888 -3344 2952 -3310
rect 2888 -3378 2892 -3344
rect 2926 -3378 2952 -3344
rect 2888 -3412 2952 -3378
rect 2888 -3446 2892 -3412
rect 2926 -3446 2952 -3412
rect 2888 -3480 2952 -3446
rect 2888 -3514 2892 -3480
rect 2926 -3514 2952 -3480
rect 2888 -3548 2952 -3514
rect 2888 -3582 2892 -3548
rect 2926 -3582 2952 -3548
rect 2888 -3610 2952 -3582
rect 4004 -2868 4090 -2810
rect 4004 -2902 4030 -2868
rect 4064 -2902 4090 -2868
rect 4004 -2936 4090 -2902
rect 4004 -2970 4030 -2936
rect 4064 -2970 4090 -2936
rect 4004 -3004 4090 -2970
rect 4004 -3038 4030 -3004
rect 4064 -3038 4090 -3004
rect 4004 -3072 4090 -3038
rect 4004 -3106 4030 -3072
rect 4064 -3106 4090 -3072
rect 4004 -3140 4090 -3106
rect 4004 -3174 4030 -3140
rect 4064 -3174 4090 -3140
rect 4004 -3208 4090 -3174
rect 4004 -3242 4030 -3208
rect 4064 -3242 4090 -3208
rect 4004 -3276 4090 -3242
rect 4004 -3310 4030 -3276
rect 4064 -3310 4090 -3276
rect 4004 -3344 4090 -3310
rect 4004 -3378 4030 -3344
rect 4064 -3378 4090 -3344
rect 4004 -3412 4090 -3378
rect 4004 -3446 4030 -3412
rect 4064 -3446 4090 -3412
rect 4004 -3480 4090 -3446
rect 4004 -3514 4030 -3480
rect 4064 -3514 4090 -3480
rect 4004 -3548 4090 -3514
rect 4004 -3582 4030 -3548
rect 4064 -3582 4090 -3548
rect 4004 -3610 4090 -3582
<< psubdiffcont >>
rect 570 -4338 650 -4166
rect 570 -4682 650 -4510
rect 570 -5026 650 -4854
rect 570 -5370 650 -5198
rect 570 -5714 650 -5542
rect 570 -6058 650 -5886
rect 570 -6402 650 -6230
rect 570 -6746 650 -6574
rect 570 -7090 650 -6918
rect 570 -7434 650 -7262
rect 570 -7778 650 -7606
rect 1176 -4338 1256 -4166
rect 1176 -4682 1256 -4510
rect 1176 -5026 1256 -4854
rect 1176 -5370 1256 -5198
rect 1176 -5714 1256 -5542
rect 1176 -6058 1256 -5886
rect 1176 -6402 1256 -6230
rect 1176 -6746 1256 -6574
rect 1176 -7090 1256 -6918
rect 1176 -7434 1256 -7262
rect 1176 -7778 1256 -7606
rect 1782 -4336 1862 -4164
rect 1782 -4680 1862 -4508
rect 1782 -5024 1862 -4852
rect 1782 -5368 1862 -5196
rect 1782 -5712 1862 -5540
rect 1782 -6056 1862 -5884
rect 1782 -6400 1862 -6228
rect 1782 -6744 1862 -6572
rect 1782 -7088 1862 -6916
rect 1782 -7432 1862 -7260
rect 1782 -7776 1862 -7604
rect 2388 -4336 2468 -4164
rect 2388 -4680 2468 -4508
rect 2388 -5024 2468 -4852
rect 2388 -5368 2468 -5196
rect 2388 -5712 2468 -5540
rect 2388 -6056 2468 -5884
rect 2388 -6400 2468 -6228
rect 2388 -6744 2468 -6572
rect 2388 -7088 2468 -6916
rect 2388 -7432 2468 -7260
rect 2388 -7776 2468 -7604
rect 2994 -4336 3074 -4164
rect 2994 -4680 3074 -4508
rect 2994 -5024 3074 -4852
rect 2994 -5368 3074 -5196
rect 2994 -5712 3074 -5540
rect 2994 -6056 3074 -5884
rect 2994 -6400 3074 -6228
rect 2994 -6744 3074 -6572
rect 2994 -7088 3074 -6916
rect 2994 -7432 3074 -7260
rect 2994 -7776 3074 -7604
rect 3600 -4336 3680 -4164
rect 3600 -4680 3680 -4508
rect 3600 -5024 3680 -4852
rect 3600 -5368 3680 -5196
rect 3600 -5712 3680 -5540
rect 3600 -6056 3680 -5884
rect 3600 -6400 3680 -6228
rect 3600 -6744 3680 -6572
rect 3600 -7088 3680 -6916
rect 3600 -7432 3680 -7260
rect 3600 -7776 3680 -7604
rect 4206 -4336 4286 -4164
rect 4206 -4680 4286 -4508
rect 4206 -5024 4286 -4852
rect 4206 -5368 4286 -5196
rect 4206 -5712 4286 -5540
rect 4206 -6056 4286 -5884
rect 4206 -6400 4286 -6228
rect 4206 -6744 4286 -6572
rect 4206 -7088 4286 -6916
rect 4206 -7432 4286 -7260
rect 4206 -7776 4286 -7604
rect 4812 -4336 4892 -4164
rect 4812 -4680 4892 -4508
rect 4812 -5024 4892 -4852
rect 4812 -5368 4892 -5196
rect 4812 -5712 4892 -5540
rect 4812 -6056 4892 -5884
rect 4812 -6400 4892 -6228
rect 4812 -6744 4892 -6572
rect 4812 -7088 4892 -6916
rect 4812 -7432 4892 -7260
rect 4812 -7776 4892 -7604
rect 5418 -4336 5498 -4164
rect 5418 -4680 5498 -4508
rect 5418 -5024 5498 -4852
rect 5418 -5368 5498 -5196
rect 5418 -5712 5498 -5540
rect 5418 -6056 5498 -5884
rect 5418 -6400 5498 -6228
rect 5418 -6744 5498 -6572
rect 5418 -7088 5498 -6916
rect 5418 -7432 5498 -7260
rect 5418 -7776 5498 -7604
rect 6024 -4336 6104 -4164
rect 6024 -4680 6104 -4508
rect 6024 -5024 6104 -4852
rect 6024 -5368 6104 -5196
rect 6024 -5712 6104 -5540
rect 6024 -6056 6104 -5884
rect 6024 -6400 6104 -6228
rect 6024 -6744 6104 -6572
rect 6024 -7088 6104 -6916
rect 6024 -7432 6104 -7260
rect 6024 -7776 6104 -7604
<< nsubdiffcont >>
rect 3498 -790 3532 -756
rect 3498 -858 3532 -824
rect 3498 -926 3532 -892
rect 3498 -994 3532 -960
rect 3498 -1062 3532 -1028
rect 3498 -1130 3532 -1096
rect 3498 -1198 3532 -1164
rect 3498 -1266 3532 -1232
rect 3498 -1334 3532 -1300
rect 3498 -1402 3532 -1368
rect 3498 -1470 3532 -1436
rect 3498 -1538 3532 -1504
rect 3498 -1606 3532 -1572
rect 3498 -1674 3532 -1640
rect 3498 -1742 3532 -1708
rect 3498 -1810 3532 -1776
rect 3498 -1878 3532 -1844
rect 3498 -1946 3532 -1912
rect 3498 -2014 3532 -1980
rect 3498 -2082 3532 -2048
rect 3498 -2150 3532 -2116
rect 3498 -2218 3532 -2184
rect 3498 -2286 3532 -2252
rect 4562 -790 4596 -756
rect 4562 -858 4596 -824
rect 4562 -926 4596 -892
rect 4562 -994 4596 -960
rect 4562 -1062 4596 -1028
rect 4562 -1130 4596 -1096
rect 4562 -1198 4596 -1164
rect 4562 -1266 4596 -1232
rect 4562 -1334 4596 -1300
rect 4562 -1402 4596 -1368
rect 4562 -1470 4596 -1436
rect 4562 -1538 4596 -1504
rect 4562 -1606 4596 -1572
rect 4562 -1674 4596 -1640
rect 4562 -1742 4596 -1708
rect 4562 -1810 4596 -1776
rect 4562 -1878 4596 -1844
rect 4562 -1946 4596 -1912
rect 4562 -2014 4596 -1980
rect 4562 -2082 4596 -2048
rect 4562 -2150 4596 -2116
rect 4562 -2218 4596 -2184
rect 4562 -2286 4596 -2252
rect 2892 -2902 2926 -2868
rect 2892 -2970 2926 -2936
rect 2892 -3038 2926 -3004
rect 2892 -3106 2926 -3072
rect 2892 -3174 2926 -3140
rect 2892 -3242 2926 -3208
rect 2892 -3310 2926 -3276
rect 2892 -3378 2926 -3344
rect 2892 -3446 2926 -3412
rect 2892 -3514 2926 -3480
rect 2892 -3582 2926 -3548
rect 4030 -2902 4064 -2868
rect 4030 -2970 4064 -2936
rect 4030 -3038 4064 -3004
rect 4030 -3106 4064 -3072
rect 4030 -3174 4064 -3140
rect 4030 -3242 4064 -3208
rect 4030 -3310 4064 -3276
rect 4030 -3378 4064 -3344
rect 4030 -3446 4064 -3412
rect 4030 -3514 4064 -3480
rect 4030 -3582 4064 -3548
<< locali >>
rect 3498 -726 3532 -710
rect 3498 -2318 3532 -2302
rect 4562 -726 4596 -710
rect 4562 -2318 4596 -2302
rect 2892 -2822 2926 -2806
rect 2892 -3614 2926 -3598
rect 4030 -2852 4064 -2806
rect 4030 -3614 4064 -3588
rect 570 -4166 650 -4150
rect 570 -7834 650 -7778
rect 1176 -4166 1256 -4150
rect 1176 -7834 1256 -7778
rect 1782 -4164 1862 -4148
rect 1782 -7832 1862 -7776
rect 2388 -4164 2468 -4148
rect 2388 -7832 2468 -7776
rect 2994 -4164 3074 -4148
rect 2994 -7832 3074 -7776
rect 3600 -4164 3680 -4148
rect 3600 -7832 3680 -7776
rect 4206 -4164 4286 -4148
rect 4206 -7832 4286 -7776
rect 4812 -4164 4892 -4148
rect 4812 -7832 4892 -7776
rect 5418 -4164 5498 -4148
rect 5418 -7832 5498 -7776
rect 6024 -4164 6104 -4148
rect 6024 -7832 6104 -7776
<< viali >>
rect 3498 -756 3532 -726
rect 3498 -790 3532 -756
rect 3498 -824 3532 -790
rect 3498 -858 3532 -824
rect 3498 -892 3532 -858
rect 3498 -926 3532 -892
rect 3498 -960 3532 -926
rect 3498 -994 3532 -960
rect 3498 -1028 3532 -994
rect 3498 -1062 3532 -1028
rect 3498 -1096 3532 -1062
rect 3498 -1130 3532 -1096
rect 3498 -1164 3532 -1130
rect 3498 -1198 3532 -1164
rect 3498 -1232 3532 -1198
rect 3498 -1266 3532 -1232
rect 3498 -1300 3532 -1266
rect 3498 -1334 3532 -1300
rect 3498 -1368 3532 -1334
rect 3498 -1402 3532 -1368
rect 3498 -1436 3532 -1402
rect 3498 -1470 3532 -1436
rect 3498 -1504 3532 -1470
rect 3498 -1538 3532 -1504
rect 3498 -1572 3532 -1538
rect 3498 -1606 3532 -1572
rect 3498 -1640 3532 -1606
rect 3498 -1674 3532 -1640
rect 3498 -1708 3532 -1674
rect 3498 -1742 3532 -1708
rect 3498 -1776 3532 -1742
rect 3498 -1810 3532 -1776
rect 3498 -1844 3532 -1810
rect 3498 -1878 3532 -1844
rect 3498 -1912 3532 -1878
rect 3498 -1946 3532 -1912
rect 3498 -1980 3532 -1946
rect 3498 -2014 3532 -1980
rect 3498 -2048 3532 -2014
rect 3498 -2082 3532 -2048
rect 3498 -2116 3532 -2082
rect 3498 -2150 3532 -2116
rect 3498 -2184 3532 -2150
rect 3498 -2218 3532 -2184
rect 3498 -2252 3532 -2218
rect 3498 -2286 3532 -2252
rect 3498 -2302 3532 -2286
rect 4562 -756 4596 -726
rect 4562 -790 4596 -756
rect 4562 -824 4596 -790
rect 4562 -858 4596 -824
rect 4562 -892 4596 -858
rect 4562 -926 4596 -892
rect 4562 -960 4596 -926
rect 4562 -994 4596 -960
rect 4562 -1028 4596 -994
rect 4562 -1062 4596 -1028
rect 4562 -1096 4596 -1062
rect 4562 -1130 4596 -1096
rect 4562 -1164 4596 -1130
rect 4562 -1198 4596 -1164
rect 4562 -1232 4596 -1198
rect 4562 -1266 4596 -1232
rect 4562 -1300 4596 -1266
rect 4562 -1334 4596 -1300
rect 4562 -1368 4596 -1334
rect 4562 -1402 4596 -1368
rect 4562 -1436 4596 -1402
rect 4562 -1470 4596 -1436
rect 4562 -1504 4596 -1470
rect 4562 -1538 4596 -1504
rect 4562 -1572 4596 -1538
rect 4562 -1606 4596 -1572
rect 4562 -1640 4596 -1606
rect 4562 -1674 4596 -1640
rect 4562 -1708 4596 -1674
rect 4562 -1742 4596 -1708
rect 4562 -1776 4596 -1742
rect 4562 -1810 4596 -1776
rect 4562 -1844 4596 -1810
rect 4562 -1878 4596 -1844
rect 4562 -1912 4596 -1878
rect 4562 -1946 4596 -1912
rect 4562 -1980 4596 -1946
rect 4562 -2014 4596 -1980
rect 4562 -2048 4596 -2014
rect 4562 -2082 4596 -2048
rect 4562 -2116 4596 -2082
rect 4562 -2150 4596 -2116
rect 4562 -2184 4596 -2150
rect 4562 -2218 4596 -2184
rect 4562 -2252 4596 -2218
rect 4562 -2286 4596 -2252
rect 4562 -2302 4596 -2286
rect 2892 -2868 2926 -2822
rect 2892 -2902 2926 -2868
rect 2892 -2936 2926 -2902
rect 2892 -2970 2926 -2936
rect 2892 -3004 2926 -2970
rect 2892 -3038 2926 -3004
rect 2892 -3072 2926 -3038
rect 2892 -3106 2926 -3072
rect 2892 -3140 2926 -3106
rect 2892 -3174 2926 -3140
rect 2892 -3208 2926 -3174
rect 2892 -3242 2926 -3208
rect 2892 -3276 2926 -3242
rect 2892 -3310 2926 -3276
rect 2892 -3344 2926 -3310
rect 2892 -3378 2926 -3344
rect 2892 -3412 2926 -3378
rect 2892 -3446 2926 -3412
rect 2892 -3480 2926 -3446
rect 2892 -3514 2926 -3480
rect 2892 -3548 2926 -3514
rect 2892 -3582 2926 -3548
rect 2892 -3598 2926 -3582
rect 4030 -2868 4064 -2852
rect 4030 -2902 4064 -2868
rect 4030 -2936 4064 -2902
rect 4030 -2970 4064 -2936
rect 4030 -3004 4064 -2970
rect 4030 -3038 4064 -3004
rect 4030 -3072 4064 -3038
rect 4030 -3106 4064 -3072
rect 4030 -3140 4064 -3106
rect 4030 -3174 4064 -3140
rect 4030 -3208 4064 -3174
rect 4030 -3242 4064 -3208
rect 4030 -3276 4064 -3242
rect 4030 -3310 4064 -3276
rect 4030 -3344 4064 -3310
rect 4030 -3378 4064 -3344
rect 4030 -3412 4064 -3378
rect 4030 -3446 4064 -3412
rect 4030 -3480 4064 -3446
rect 4030 -3514 4064 -3480
rect 4030 -3548 4064 -3514
rect 4030 -3582 4064 -3548
rect 4030 -3588 4064 -3582
rect 570 -4338 650 -4166
rect 570 -4510 650 -4338
rect 570 -4682 650 -4510
rect 570 -4854 650 -4682
rect 570 -5026 650 -4854
rect 570 -5198 650 -5026
rect 570 -5370 650 -5198
rect 570 -5542 650 -5370
rect 570 -5714 650 -5542
rect 570 -5886 650 -5714
rect 570 -6058 650 -5886
rect 570 -6230 650 -6058
rect 570 -6402 650 -6230
rect 570 -6574 650 -6402
rect 570 -6746 650 -6574
rect 570 -6918 650 -6746
rect 570 -7090 650 -6918
rect 570 -7262 650 -7090
rect 570 -7434 650 -7262
rect 570 -7606 650 -7434
rect 570 -7778 650 -7606
rect 1176 -4338 1256 -4166
rect 1176 -4510 1256 -4338
rect 1176 -4682 1256 -4510
rect 1176 -4854 1256 -4682
rect 1176 -5026 1256 -4854
rect 1176 -5198 1256 -5026
rect 1176 -5370 1256 -5198
rect 1176 -5542 1256 -5370
rect 1176 -5714 1256 -5542
rect 1176 -5886 1256 -5714
rect 1176 -6058 1256 -5886
rect 1176 -6230 1256 -6058
rect 1176 -6402 1256 -6230
rect 1176 -6574 1256 -6402
rect 1176 -6746 1256 -6574
rect 1176 -6918 1256 -6746
rect 1176 -7090 1256 -6918
rect 1176 -7262 1256 -7090
rect 1176 -7434 1256 -7262
rect 1176 -7606 1256 -7434
rect 1176 -7778 1256 -7606
rect 1782 -4336 1862 -4164
rect 1782 -4508 1862 -4336
rect 1782 -4680 1862 -4508
rect 1782 -4852 1862 -4680
rect 1782 -5024 1862 -4852
rect 1782 -5196 1862 -5024
rect 1782 -5368 1862 -5196
rect 1782 -5540 1862 -5368
rect 1782 -5712 1862 -5540
rect 1782 -5884 1862 -5712
rect 1782 -6056 1862 -5884
rect 1782 -6228 1862 -6056
rect 1782 -6400 1862 -6228
rect 1782 -6572 1862 -6400
rect 1782 -6744 1862 -6572
rect 1782 -6916 1862 -6744
rect 1782 -7088 1862 -6916
rect 1782 -7260 1862 -7088
rect 1782 -7432 1862 -7260
rect 1782 -7604 1862 -7432
rect 1782 -7776 1862 -7604
rect 2388 -4336 2468 -4164
rect 2388 -4508 2468 -4336
rect 2388 -4680 2468 -4508
rect 2388 -4852 2468 -4680
rect 2388 -5024 2468 -4852
rect 2388 -5196 2468 -5024
rect 2388 -5368 2468 -5196
rect 2388 -5540 2468 -5368
rect 2388 -5712 2468 -5540
rect 2388 -5884 2468 -5712
rect 2388 -6056 2468 -5884
rect 2388 -6228 2468 -6056
rect 2388 -6400 2468 -6228
rect 2388 -6572 2468 -6400
rect 2388 -6744 2468 -6572
rect 2388 -6916 2468 -6744
rect 2388 -7088 2468 -6916
rect 2388 -7260 2468 -7088
rect 2388 -7432 2468 -7260
rect 2388 -7604 2468 -7432
rect 2388 -7776 2468 -7604
rect 2994 -4336 3074 -4164
rect 2994 -4508 3074 -4336
rect 2994 -4680 3074 -4508
rect 2994 -4852 3074 -4680
rect 2994 -5024 3074 -4852
rect 2994 -5196 3074 -5024
rect 2994 -5368 3074 -5196
rect 2994 -5540 3074 -5368
rect 2994 -5712 3074 -5540
rect 2994 -5884 3074 -5712
rect 2994 -6056 3074 -5884
rect 2994 -6228 3074 -6056
rect 2994 -6400 3074 -6228
rect 2994 -6572 3074 -6400
rect 2994 -6744 3074 -6572
rect 2994 -6916 3074 -6744
rect 2994 -7088 3074 -6916
rect 2994 -7260 3074 -7088
rect 2994 -7432 3074 -7260
rect 2994 -7604 3074 -7432
rect 2994 -7776 3074 -7604
rect 3600 -4336 3680 -4164
rect 3600 -4508 3680 -4336
rect 3600 -4680 3680 -4508
rect 3600 -4852 3680 -4680
rect 3600 -5024 3680 -4852
rect 3600 -5196 3680 -5024
rect 3600 -5368 3680 -5196
rect 3600 -5540 3680 -5368
rect 3600 -5712 3680 -5540
rect 3600 -5884 3680 -5712
rect 3600 -6056 3680 -5884
rect 3600 -6228 3680 -6056
rect 3600 -6400 3680 -6228
rect 3600 -6572 3680 -6400
rect 3600 -6744 3680 -6572
rect 3600 -6916 3680 -6744
rect 3600 -7088 3680 -6916
rect 3600 -7260 3680 -7088
rect 3600 -7432 3680 -7260
rect 3600 -7604 3680 -7432
rect 3600 -7776 3680 -7604
rect 4206 -4336 4286 -4164
rect 4206 -4508 4286 -4336
rect 4206 -4680 4286 -4508
rect 4206 -4852 4286 -4680
rect 4206 -5024 4286 -4852
rect 4206 -5196 4286 -5024
rect 4206 -5368 4286 -5196
rect 4206 -5540 4286 -5368
rect 4206 -5712 4286 -5540
rect 4206 -5884 4286 -5712
rect 4206 -6056 4286 -5884
rect 4206 -6228 4286 -6056
rect 4206 -6400 4286 -6228
rect 4206 -6572 4286 -6400
rect 4206 -6744 4286 -6572
rect 4206 -6916 4286 -6744
rect 4206 -7088 4286 -6916
rect 4206 -7260 4286 -7088
rect 4206 -7432 4286 -7260
rect 4206 -7604 4286 -7432
rect 4206 -7776 4286 -7604
rect 4812 -4336 4892 -4164
rect 4812 -4508 4892 -4336
rect 4812 -4680 4892 -4508
rect 4812 -4852 4892 -4680
rect 4812 -5024 4892 -4852
rect 4812 -5196 4892 -5024
rect 4812 -5368 4892 -5196
rect 4812 -5540 4892 -5368
rect 4812 -5712 4892 -5540
rect 4812 -5884 4892 -5712
rect 4812 -6056 4892 -5884
rect 4812 -6228 4892 -6056
rect 4812 -6400 4892 -6228
rect 4812 -6572 4892 -6400
rect 4812 -6744 4892 -6572
rect 4812 -6916 4892 -6744
rect 4812 -7088 4892 -6916
rect 4812 -7260 4892 -7088
rect 4812 -7432 4892 -7260
rect 4812 -7604 4892 -7432
rect 4812 -7776 4892 -7604
rect 5418 -4336 5498 -4164
rect 5418 -4508 5498 -4336
rect 5418 -4680 5498 -4508
rect 5418 -4852 5498 -4680
rect 5418 -5024 5498 -4852
rect 5418 -5196 5498 -5024
rect 5418 -5368 5498 -5196
rect 5418 -5540 5498 -5368
rect 5418 -5712 5498 -5540
rect 5418 -5884 5498 -5712
rect 5418 -6056 5498 -5884
rect 5418 -6228 5498 -6056
rect 5418 -6400 5498 -6228
rect 5418 -6572 5498 -6400
rect 5418 -6744 5498 -6572
rect 5418 -6916 5498 -6744
rect 5418 -7088 5498 -6916
rect 5418 -7260 5498 -7088
rect 5418 -7432 5498 -7260
rect 5418 -7604 5498 -7432
rect 5418 -7776 5498 -7604
rect 6024 -4336 6104 -4164
rect 6024 -4508 6104 -4336
rect 6024 -4680 6104 -4508
rect 6024 -4852 6104 -4680
rect 6024 -5024 6104 -4852
rect 6024 -5196 6104 -5024
rect 6024 -5368 6104 -5196
rect 6024 -5540 6104 -5368
rect 6024 -5712 6104 -5540
rect 6024 -5884 6104 -5712
rect 6024 -6056 6104 -5884
rect 6024 -6228 6104 -6056
rect 6024 -6400 6104 -6228
rect 6024 -6572 6104 -6400
rect 6024 -6744 6104 -6572
rect 6024 -6916 6104 -6744
rect 6024 -7088 6104 -6916
rect 6024 -7260 6104 -7088
rect 6024 -7432 6104 -7260
rect 6024 -7604 6104 -7432
rect 6024 -7776 6104 -7604
<< metal1 >>
rect 2814 -104 2870 -98
rect 2814 -454 2816 -104
rect 2868 -454 2870 -104
rect 4 -2330 228 -1140
rect 4 -2426 12 -2330
rect 220 -2426 228 -2330
rect 4 -2434 228 -2426
rect 4 -2652 228 -2644
rect 4 -3726 10 -2652
rect 220 -3626 228 -2652
rect 2814 -2810 2870 -454
rect 3458 -104 3572 -98
rect 3458 -454 3466 -104
rect 3564 -454 3572 -104
rect 3458 -726 3572 -454
rect 4488 -104 4732 -96
rect 4488 -454 4496 -104
rect 4726 -454 4732 -104
rect 4488 -614 4732 -454
rect 4488 -714 4602 -614
rect 4528 -726 4602 -714
rect 2954 -778 3012 -768
rect 2954 -2268 3012 -2258
rect 3464 -2302 3498 -726
rect 3532 -2302 3566 -726
rect 4018 -778 4076 -768
rect 4018 -2268 4076 -2258
rect 3464 -2314 3566 -2302
rect 4528 -2302 4562 -726
rect 4596 -2302 4602 -726
rect 4528 -2314 4602 -2302
rect 3022 -2406 3028 -2350
rect 3396 -2406 3402 -2350
rect 3628 -2406 3634 -2350
rect 4002 -2406 4008 -2350
rect 4086 -2406 4092 -2350
rect 4460 -2406 4466 -2350
rect 3756 -2608 3868 -2544
rect 3756 -2728 3764 -2608
rect 3860 -2728 3868 -2608
rect 2814 -2822 2932 -2810
rect 2814 -3598 2892 -2822
rect 2926 -3598 2932 -2822
rect 2966 -2882 3026 -2870
rect 2966 -3568 3026 -3556
rect 2814 -3610 2932 -3598
rect 3088 -3610 3288 -2810
rect 3756 -3610 3868 -2728
rect 4226 -2608 4338 -2544
rect 4226 -2728 4234 -2608
rect 4330 -2728 4338 -2608
rect 3944 -2886 3996 -2810
rect 3944 -3610 3996 -3554
rect 4024 -2852 4070 -2810
rect 4024 -3588 4030 -2852
rect 4064 -3588 4070 -2852
rect 4024 -3610 4070 -3588
rect 4098 -2886 4150 -2810
rect 4098 -3610 4150 -3554
rect 4226 -3610 4338 -2728
rect 222 -3726 228 -3626
rect 3012 -3644 3082 -3638
rect 3012 -3706 3082 -3700
rect 4 -3732 228 -3726
rect 6 -3804 230 -3794
rect 6 -3896 16 -3804
rect 220 -3896 230 -3804
rect 6 -5088 230 -3896
rect 3176 -3804 3288 -3610
rect 3874 -3644 3944 -3638
rect 3874 -3706 3944 -3700
rect 3176 -3896 3186 -3804
rect 3278 -3896 3288 -3804
rect 4030 -3804 4064 -3610
rect 4150 -3644 4220 -3638
rect 4150 -3706 4220 -3700
rect 4676 -3804 4732 -614
rect 6388 -2552 6838 -1412
rect 6388 -2760 6396 -2552
rect 6830 -2760 6838 -2552
rect 6388 -2768 6838 -2760
rect 4030 -3808 4106 -3804
rect 4030 -3860 4036 -3808
rect 4100 -3860 4106 -3808
rect 4618 -3808 4732 -3804
rect 4618 -3860 4628 -3808
rect 4726 -3860 4732 -3808
rect 774 -3968 1056 -3962
rect 774 -4124 788 -3968
rect 1046 -4124 1056 -3968
rect 3176 -3968 3288 -3896
rect 3176 -4124 3182 -3968
rect 3282 -4124 3288 -3968
rect 564 -4166 656 -4150
rect 774 -4164 1056 -4124
rect 564 -7778 570 -4166
rect 650 -7778 656 -4166
rect 1170 -4166 1262 -4150
rect 1776 -4164 1868 -4148
rect 564 -7926 656 -7778
rect 790 -7420 1040 -7414
rect 790 -7822 1040 -7816
rect 1170 -7778 1176 -4166
rect 1256 -7778 1262 -4166
rect 1396 -4170 1646 -4164
rect 1396 -4572 1646 -4566
rect 564 -8358 572 -7926
rect 648 -8358 656 -7926
rect 564 -8366 656 -8358
rect 1170 -7926 1262 -7778
rect 1396 -7420 1646 -7414
rect 1396 -7822 1646 -7816
rect 1776 -7776 1782 -4164
rect 1862 -7776 1868 -4164
rect 2002 -4168 2252 -4162
rect 2002 -4570 2252 -4564
rect 2382 -4164 2474 -4148
rect 1170 -8358 1178 -7926
rect 1254 -8358 1262 -7926
rect 1170 -8366 1262 -8358
rect 1776 -7926 1868 -7776
rect 2002 -7418 2252 -7412
rect 2002 -7820 2252 -7814
rect 2382 -7776 2388 -4164
rect 2468 -7776 2474 -4164
rect 2608 -4168 2858 -4162
rect 2608 -4570 2858 -4564
rect 2988 -4164 3080 -4148
rect 1776 -8358 1784 -7926
rect 1860 -8358 1868 -7926
rect 1776 -8366 1868 -8358
rect 2382 -7926 2474 -7776
rect 2608 -7418 2858 -7412
rect 2608 -7820 2858 -7814
rect 2988 -7776 2994 -4164
rect 3074 -7776 3080 -4164
rect 3214 -4168 3464 -4162
rect 3214 -4570 3464 -4564
rect 3594 -4164 3686 -4148
rect 2382 -8358 2390 -7926
rect 2466 -8358 2474 -7926
rect 2382 -8366 2474 -8358
rect 2988 -7926 3080 -7776
rect 3214 -7418 3464 -7412
rect 3214 -7820 3464 -7814
rect 3594 -7776 3600 -4164
rect 3680 -7776 3686 -4164
rect 3820 -4168 4070 -4162
rect 3820 -4570 4070 -4564
rect 4200 -4164 4292 -4148
rect 2988 -8358 2996 -7926
rect 3072 -8358 3080 -7926
rect 2988 -8366 3080 -8358
rect 3594 -7926 3686 -7776
rect 3820 -7418 4070 -7412
rect 3820 -7820 4070 -7814
rect 4200 -7776 4206 -4164
rect 4286 -7776 4292 -4164
rect 4426 -4168 4676 -4162
rect 4426 -4570 4676 -4564
rect 4806 -4164 4898 -4148
rect 3594 -8358 3602 -7926
rect 3678 -8358 3686 -7926
rect 3594 -8366 3686 -8358
rect 4200 -7926 4292 -7776
rect 4426 -7418 4676 -7412
rect 4426 -7820 4676 -7814
rect 4806 -7776 4812 -4164
rect 4892 -7776 4898 -4164
rect 5032 -4168 5282 -4162
rect 5032 -4570 5282 -4564
rect 5412 -4164 5504 -4148
rect 4200 -8358 4208 -7926
rect 4284 -8358 4292 -7926
rect 4200 -8366 4292 -8358
rect 4806 -7926 4898 -7776
rect 5032 -7418 5282 -7412
rect 5032 -7820 5282 -7814
rect 5412 -7776 5418 -4164
rect 5498 -7776 5504 -4164
rect 5638 -4168 5888 -4162
rect 5638 -4570 5888 -4564
rect 6018 -4164 6110 -4148
rect 4806 -8358 4814 -7926
rect 4890 -8358 4898 -7926
rect 4806 -8366 4898 -8358
rect 5412 -7926 5504 -7776
rect 5638 -7418 5888 -7412
rect 5638 -7820 5888 -7814
rect 6018 -7776 6024 -4164
rect 6104 -7776 6110 -4164
rect 6244 -4168 6494 -4162
rect 6244 -4570 6494 -4564
rect 6600 -4168 6768 -4160
rect 6600 -4562 6608 -4168
rect 6760 -4562 6768 -4168
rect 5412 -8358 5420 -7926
rect 5496 -8358 5504 -7926
rect 5412 -8366 5504 -8358
rect 6018 -7926 6110 -7776
rect 6244 -7418 6494 -7412
rect 6244 -7820 6494 -7814
rect 6018 -8358 6026 -7926
rect 6102 -8358 6110 -7926
rect 6018 -8366 6110 -8358
rect 6600 -7918 6768 -4562
rect 6600 -7926 6776 -7918
rect 6600 -8358 6608 -7926
rect 6764 -8358 6776 -7926
rect 6600 -8366 6776 -8358
<< via1 >>
rect 2816 -454 2868 -104
rect 12 -2426 220 -2330
rect 10 -3626 220 -2652
rect 3466 -454 3564 -104
rect 4496 -454 4726 -104
rect 2954 -2258 3012 -778
rect 4018 -2258 4076 -778
rect 3028 -2406 3396 -2350
rect 3634 -2406 4002 -2350
rect 4092 -2406 4460 -2350
rect 3764 -2728 3860 -2608
rect 2966 -3556 3026 -2882
rect 4234 -2728 4330 -2608
rect 3944 -3554 3996 -2886
rect 4098 -3554 4150 -2886
rect 10 -3726 222 -3626
rect 3012 -3700 3082 -3644
rect 16 -3896 220 -3804
rect 3874 -3700 3944 -3644
rect 3186 -3896 3278 -3804
rect 4150 -3700 4220 -3644
rect 6396 -2760 6830 -2552
rect 4036 -3860 4100 -3808
rect 4628 -3860 4726 -3808
rect 788 -4124 1046 -3968
rect 3182 -4124 3282 -3968
rect 790 -7816 1040 -7420
rect 1396 -4566 1646 -4170
rect 572 -8358 648 -7926
rect 1396 -7816 1646 -7420
rect 2002 -4564 2252 -4168
rect 1178 -8358 1254 -7926
rect 2002 -7814 2252 -7418
rect 2608 -4564 2858 -4168
rect 1784 -8358 1860 -7926
rect 2608 -7814 2858 -7418
rect 3214 -4564 3464 -4168
rect 2390 -8358 2466 -7926
rect 3214 -7814 3464 -7418
rect 3820 -4564 4070 -4168
rect 2996 -8358 3072 -7926
rect 3820 -7814 4070 -7418
rect 4426 -4564 4676 -4168
rect 3602 -8358 3678 -7926
rect 4426 -7814 4676 -7418
rect 5032 -4564 5282 -4168
rect 4208 -8358 4284 -7926
rect 5032 -7814 5282 -7418
rect 5638 -4564 5888 -4168
rect 4814 -8358 4890 -7926
rect 5638 -7814 5888 -7418
rect 6244 -4564 6494 -4168
rect 6608 -4562 6760 -4168
rect 5420 -8358 5496 -7926
rect 6244 -7814 6494 -7418
rect 6026 -8358 6102 -7926
rect 6608 -8358 6764 -7926
<< metal2 >>
rect 4 -104 6836 -32
rect 4 -454 2816 -104
rect 2868 -454 3466 -104
rect 3564 -454 4496 -104
rect 4726 -454 6836 -104
rect 4 -480 6836 -454
rect 2954 -778 3012 -768
rect 2954 -2268 3012 -2258
rect 4018 -778 4076 -768
rect 4018 -2268 4076 -2258
rect 4 -2330 4480 -2322
rect 4 -2426 12 -2330
rect 220 -2332 4480 -2330
rect 220 -2424 2654 -2332
rect 2762 -2350 4480 -2332
rect 2762 -2406 3028 -2350
rect 3396 -2406 3634 -2350
rect 4002 -2406 4092 -2350
rect 4460 -2406 4480 -2350
rect 2762 -2424 4480 -2406
rect 220 -2426 4480 -2424
rect 4 -2434 4480 -2426
rect 3756 -2552 6838 -2544
rect 3756 -2608 6396 -2552
rect 4 -2652 228 -2644
rect 4 -3726 10 -2652
rect 220 -3620 228 -2652
rect 3756 -2728 3764 -2608
rect 3860 -2728 4234 -2608
rect 4330 -2728 6396 -2608
rect 3756 -2760 6396 -2728
rect 6830 -2760 6838 -2552
rect 3756 -2768 6838 -2760
rect 2966 -2882 3026 -2870
rect 2966 -3568 3026 -3556
rect 3944 -2886 4002 -2876
rect 3944 -3564 4002 -3554
rect 4092 -2886 4150 -2876
rect 4092 -3564 4150 -3554
rect 220 -3626 4242 -3620
rect 222 -3644 4242 -3626
rect 222 -3700 3012 -3644
rect 3082 -3700 3874 -3644
rect 3944 -3700 4150 -3644
rect 4220 -3700 4242 -3644
rect 222 -3726 4242 -3700
rect 4 -3732 4242 -3726
rect 6 -3804 230 -3794
rect 6 -3896 16 -3804
rect 220 -3896 230 -3804
rect 6 -3906 230 -3896
rect 3176 -3804 3288 -3794
rect 3176 -3896 3186 -3804
rect 3278 -3896 3288 -3804
rect 4030 -3808 4732 -3804
rect 4030 -3860 4036 -3808
rect 4100 -3860 4628 -3808
rect 4726 -3860 4732 -3808
rect 3176 -3906 3288 -3896
rect 774 -3968 3288 -3962
rect 774 -4124 788 -3968
rect 1046 -4124 3182 -3968
rect 3282 -4124 3288 -3968
rect 774 -4130 3288 -4124
rect 2856 -4162 3216 -4160
rect 4068 -4162 4428 -4160
rect 5280 -4162 5640 -4160
rect 1396 -4168 2252 -4162
rect 1396 -4170 2002 -4168
rect 1646 -4564 2002 -4170
rect 1646 -4566 2252 -4564
rect 1396 -4572 2252 -4566
rect 2608 -4168 3464 -4162
rect 2858 -4564 3214 -4168
rect 2608 -4570 3464 -4564
rect 3820 -4168 4676 -4162
rect 4070 -4564 4426 -4168
rect 3820 -4570 4676 -4564
rect 5032 -4168 5888 -4162
rect 5282 -4564 5638 -4168
rect 5032 -4570 5888 -4564
rect 6244 -4168 6768 -4160
rect 6494 -4562 6608 -4168
rect 6760 -4562 6768 -4168
rect 6494 -4564 6768 -4562
rect 6244 -4570 6768 -4564
rect 2250 -7412 2610 -7410
rect 3462 -7412 3822 -7410
rect 4674 -7412 5034 -7410
rect 5886 -7412 6494 -7410
rect 790 -7420 1646 -7414
rect 1040 -7816 1396 -7420
rect 790 -7822 1646 -7816
rect 2002 -7418 2858 -7412
rect 2252 -7814 2608 -7418
rect 2002 -7820 2858 -7814
rect 3214 -7418 4070 -7412
rect 3464 -7814 3820 -7418
rect 3214 -7820 4070 -7814
rect 4426 -7418 5282 -7412
rect 4676 -7814 5032 -7418
rect 4426 -7820 5282 -7814
rect 5638 -7418 6494 -7412
rect 5888 -7814 6244 -7418
rect 5638 -7820 6494 -7814
rect 546 -7926 6836 -7918
rect 546 -8358 572 -7926
rect 648 -8358 1178 -7926
rect 1254 -8358 1784 -7926
rect 1860 -8358 2390 -7926
rect 2466 -8358 2996 -7926
rect 3072 -8358 3602 -7926
rect 3678 -8358 4208 -7926
rect 4284 -8358 4814 -7926
rect 4890 -8358 5420 -7926
rect 5496 -8358 6026 -7926
rect 6102 -8358 6608 -7926
rect 6764 -8358 6836 -7926
rect 546 -8366 6836 -8358
<< via2 >>
rect 2954 -2258 3012 -778
rect 4018 -2258 4076 -778
rect 2654 -2424 2762 -2332
rect 2966 -3556 3026 -2882
rect 3944 -3554 3996 -2886
rect 3996 -3554 4002 -2886
rect 4092 -3554 4098 -2886
rect 4098 -3554 4150 -2886
rect 16 -3896 220 -3804
rect 3186 -3896 3278 -3804
<< metal3 >>
rect 2934 -778 3054 -760
rect 2934 -2258 2954 -778
rect 3012 -2258 3054 -778
rect 2646 -2332 2770 -2322
rect 2646 -2424 2654 -2332
rect 2762 -2424 2770 -2332
rect 2646 -2434 2770 -2424
rect 2934 -2882 3054 -2258
rect 3956 -778 4136 -762
rect 3956 -2258 4018 -778
rect 4076 -2258 4136 -778
rect 3956 -2876 4136 -2258
rect 2934 -3556 2966 -2882
rect 3026 -3556 3054 -2882
rect 2934 -3568 3054 -3556
rect 3938 -2886 4156 -2876
rect 3938 -3554 3944 -2886
rect 4002 -3554 4092 -2886
rect 4150 -3554 4156 -2886
rect 3938 -3564 4156 -3554
rect 6 -3804 230 -3794
rect 6 -3896 16 -3804
rect 220 -3896 230 -3804
rect 6 -3906 230 -3896
rect 3176 -3804 3288 -3794
rect 3176 -3896 3186 -3804
rect 3278 -3896 3288 -3804
rect 3176 -3906 3288 -3896
<< via3 >>
rect 2654 -2424 2762 -2332
rect 16 -3896 220 -3804
rect 3186 -3896 3278 -3804
<< metal4 >>
rect 1566 -2332 2770 -2322
rect 1566 -2424 2654 -2332
rect 2762 -2424 2770 -2332
rect 1566 -2434 2770 -2424
rect 1566 -2520 2566 -2434
rect 1498 -3794 2554 -3790
rect 6 -3804 3288 -3794
rect 6 -3896 16 -3804
rect 220 -3896 3186 -3804
rect 3278 -3896 3288 -3804
rect 6 -3906 3288 -3896
use sky130_fd_pr__pfet_01v8_lvt_HL7PVG  M1
timestamp 1681673980
transform -1 0 3212 0 1 -1550
box -294 -864 294 898
use sky130_fd_pr__pfet_01v8_lvt_73XLH3  M2
timestamp 1680972802
transform 1 0 3047 0 1 -3246
box -129 -464 129 498
use sky130_fd_pr__pfet_01v8_lvt_HL7PVG  M31
timestamp 1681673980
transform 1 0 3818 0 1 -1550
box -294 -864 294 898
use sky130_fd_pr__pfet_01v8_lvt_HL7PVG  M32
timestamp 1681673980
transform -1 0 4276 0 1 -1550
box -294 -864 294 898
use sky130_fd_pr__pfet_01v8_lvt_73XLH3  M41
timestamp 1680972802
transform -1 0 3909 0 1 -3246
box -129 -464 129 498
use sky130_fd_pr__pfet_01v8_lvt_73XLH3  M42
timestamp 1680972802
transform 1 0 4185 0 1 -3246
box -129 -464 129 498
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  XC1
timestamp 1680255405
transform 0 1 2026 -1 0 -3120
box -686 -540 686 540
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR11
timestamp 1680448829
transform 1 0 915 0 1 -5992
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_TE7XP6  XR12
timestamp 1680449562
transform 1 0 1521 0 1 -5992
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR13
timestamp 1680448829
transform 1 0 2127 0 1 -5990
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR14
timestamp 1680448829
transform 1 0 2733 0 1 -5990
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR15
timestamp 1680448829
transform 1 0 3339 0 1 -5990
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR16
timestamp 1680448829
transform 1 0 3945 0 1 -5990
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_CW7864  XR17
timestamp 1680448829
transform 1 0 4551 0 1 -5990
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_TE7XP6  XR18
timestamp 1680449562
transform 1 0 5157 0 1 -5990
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_TE7XP6  XR19
timestamp 1680449562
transform 1 0 5763 0 1 -5990
box -143 -1842 143 1842
use sky130_fd_pr__res_xhigh_po_1p41_TE7XP6  XR20
timestamp 1680449562
transform 1 0 6369 0 1 -5990
box -143 -1842 143 1842
<< labels >>
flabel metal2 546 -8366 6836 -7918 0 FreeMono 2400 0 0 0 vss
port 1 nsew
flabel metal1 6388 -2768 6838 -1412 0 FreeMono 2400 90 0 0 iout
port 2 nsew
flabel metal1 6 -5088 230 -3794 0 FreeMono 1120 90 0 0 fb
port 5 nsew
flabel metal1 4 -2434 228 -1140 0 FreeMono 1120 90 0 0 outop
port 4 nsew
flabel metal1 4 -3732 228 -2644 0 FreeMono 1120 90 0 0 bgr
port 3 nsew
flabel metal2 4 -480 6836 -32 0 FreeMono 2400 0 0 0 vdd
port 0 nsew
<< end >>
