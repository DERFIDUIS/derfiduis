magic
tech sky130A
magscale 1 2
timestamp 1681050310
<< error_p >>
rect -31 -511 31 -505
rect -31 -545 -19 -511
rect -31 -551 31 -545
<< nwell >>
rect -129 -564 129 598
<< pmoslvt >>
rect -35 -464 35 536
<< pdiff >>
rect -93 524 -35 536
rect -93 -452 -81 524
rect -47 -452 -35 524
rect -93 -464 -35 -452
rect 35 524 93 536
rect 35 -452 47 524
rect 81 -452 93 524
rect 35 -464 93 -452
<< pdiffc >>
rect -81 -452 -47 524
rect 47 -452 81 524
<< poly >>
rect -35 536 35 562
rect -35 -511 35 -464
rect -35 -545 -19 -511
rect 19 -545 35 -511
rect -35 -561 35 -545
<< polycont >>
rect -19 -545 19 -511
<< locali >>
rect -81 524 -47 540
rect -81 -468 -47 -452
rect 47 524 81 540
rect 47 -468 81 -452
rect -35 -545 -19 -511
rect 19 -545 35 -511
<< viali >>
rect -81 -452 -47 524
rect 47 -452 81 524
rect -19 -545 19 -511
<< metal1 >>
rect -87 524 -41 536
rect -87 -452 -81 524
rect -47 -452 -41 524
rect -87 -464 -41 -452
rect 41 524 87 536
rect 41 -452 47 524
rect 81 -452 87 524
rect 41 -464 87 -452
rect -31 -511 31 -505
rect -31 -545 -19 -511
rect 19 -545 31 -511
rect -31 -551 31 -545
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 5.0 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
