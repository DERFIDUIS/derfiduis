magic
tech sky130A
magscale 1 2
timestamp 1680265380
<< error_p >>
rect -29 572 29 578
rect -29 538 -17 572
rect -29 532 29 538
rect -29 -538 29 -532
rect -29 -572 -17 -538
rect -29 -578 29 -572
<< pwell >>
rect -214 -710 214 710
<< nmoslvt >>
rect -18 -500 18 500
<< ndiff >>
rect -76 488 -18 500
rect -76 -488 -64 488
rect -30 -488 -18 488
rect -76 -500 -18 -488
rect 18 488 76 500
rect 18 -488 30 488
rect 64 -488 76 488
rect 18 -500 76 -488
<< ndiffc >>
rect -64 -488 -30 488
rect 30 -488 64 488
<< psubdiff >>
rect -178 640 -82 674
rect 82 640 178 674
rect -178 578 -144 640
rect 144 578 178 640
rect -178 -640 -144 -578
rect 144 -640 178 -578
rect -178 -674 -82 -640
rect 82 -674 178 -640
<< psubdiffcont >>
rect -82 640 82 674
rect -178 -578 -144 578
rect 144 -578 178 578
rect -82 -674 82 -640
<< poly >>
rect -33 572 33 588
rect -33 538 -17 572
rect 17 538 33 572
rect -33 522 33 538
rect -18 500 18 522
rect -18 -522 18 -500
rect -33 -538 33 -522
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect -33 -588 33 -572
<< polycont >>
rect -17 538 17 572
rect -17 -572 17 -538
<< locali >>
rect -178 640 -82 674
rect 82 640 178 674
rect -178 578 -144 640
rect 144 578 178 640
rect -33 538 -17 572
rect 17 538 33 572
rect -64 488 -30 504
rect -64 -504 -30 -488
rect 30 488 64 504
rect 30 -504 64 -488
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect -178 -640 -144 -578
rect 144 -640 178 -578
rect -178 -674 -82 -640
rect 82 -674 178 -640
<< viali >>
rect -17 538 17 572
rect -64 -488 -30 488
rect 30 -488 64 488
rect -17 -572 17 -538
<< metal1 >>
rect -29 572 29 578
rect -29 538 -17 572
rect 17 538 29 572
rect -29 532 29 538
rect -70 488 -24 500
rect -70 -488 -64 488
rect -30 -488 -24 488
rect -70 -500 -24 -488
rect 24 488 70 500
rect 24 -488 30 488
rect 64 -488 70 488
rect 24 -500 70 -488
rect -29 -538 29 -532
rect -29 -572 -17 -538
rect 17 -572 29 -538
rect -29 -578 29 -572
<< properties >>
string FIXED_BBOX -161 -657 161 657
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 5.0 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
