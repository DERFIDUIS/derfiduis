** sch_path: /home/karlajcm/Documentos/TESIS DE
*+ GRADO/WORK_IN_PROGRESS/My_xschem/For_Layout/rectifier_lvt_01v8_initial.sch
.subckt rectifier_lvt_01v8_initial vinp vinn vss out2
*.PININFO vinp:B vinn:B vss:B out2:B
M11 vinp vinn vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M21 vinn vinp vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M31 vinp vinn out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M41 vinn vinp out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M12 vinp vinn vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M13 vinp vinn vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M14 vinp vinn vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M15 vinp vinn vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M16 vinp vinn vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M22 vinn vinp vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M23 vinn vinp vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M24 vinn vinp vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M25 vinn vinp vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M26 vinn vinp vss vss sky130_fd_pr__nfet_01v8_lvt L=0.18 W=5 nf=1 m=1
M32 vinp vinn out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M33 vinp vinn out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M34 vinp vinn out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M35 vinp vinn out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M36 vinp vinn out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M42 vinn vinp out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M43 vinn vinp out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M44 vinn vinp out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M45 vinn vinp out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
M46 vinn vinp out2 out2 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=5 nf=1 m=1
.ends
.end
