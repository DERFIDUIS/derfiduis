magic
tech sky130A
magscale 1 2
timestamp 1680985943
<< error_p >>
rect -129 -498 129 464
<< nwell >>
rect -129 -498 129 464
<< pmoslvt >>
rect -35 -436 35 364
<< pdiff >>
rect -93 352 -35 364
rect -93 -424 -81 352
rect -47 -424 -35 352
rect -93 -436 -35 -424
rect 35 352 93 364
rect 35 -424 47 352
rect 81 -424 93 352
rect 35 -436 93 -424
<< pdiffc >>
rect -81 -424 -47 352
rect 47 -424 81 352
<< poly >>
rect -35 445 35 461
rect -35 411 -19 445
rect 19 411 35 445
rect -35 364 35 411
rect -35 -462 35 -436
<< polycont >>
rect -19 411 19 445
<< locali >>
rect -35 411 -19 445
rect 19 411 35 445
rect -81 352 -47 368
rect -81 -440 -47 -424
rect 47 352 81 368
rect 47 -440 81 -424
<< viali >>
rect -19 411 19 445
rect -81 -424 -47 352
rect 47 -424 81 352
<< metal1 >>
rect -31 445 31 451
rect -31 411 -19 445
rect 19 411 31 445
rect -31 405 31 411
rect -87 352 -41 364
rect -87 -424 -81 352
rect -47 -424 -41 352
rect -87 -436 -41 -424
rect 41 352 87 364
rect 41 -424 47 352
rect 81 -424 87 352
rect 41 -436 87 -424
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 4.0 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
