magic
tech sky130A
magscale 1 2
timestamp 1680254034
<< nwell >>
rect -294 -1300 294 1300
<< pmoslvt >>
rect -200 -1200 200 1200
<< pdiff >>
rect -258 1188 -200 1200
rect -258 -1188 -246 1188
rect -212 -1188 -200 1188
rect -258 -1200 -200 -1188
rect 200 1188 258 1200
rect 200 -1188 212 1188
rect 246 -1188 258 1188
rect 200 -1200 258 -1188
<< pdiffc >>
rect -246 -1188 -212 1188
rect 212 -1188 246 1188
<< poly >>
rect -200 1281 200 1297
rect -200 1247 -184 1281
rect 184 1247 200 1281
rect -200 1200 200 1247
rect -200 -1247 200 -1200
rect -200 -1281 -184 -1247
rect 184 -1281 200 -1247
rect -200 -1297 200 -1281
<< polycont >>
rect -184 1247 184 1281
rect -184 -1281 184 -1247
<< locali >>
rect -200 1247 -184 1281
rect 184 1247 200 1281
rect -246 1188 -212 1204
rect -246 -1204 -212 -1188
rect 212 1188 246 1204
rect 212 -1204 246 -1188
rect -200 -1281 -184 -1247
rect 184 -1281 200 -1247
<< viali >>
rect -184 1247 184 1281
rect -246 -1188 -212 1188
rect 212 -1188 246 1188
rect -184 -1281 184 -1247
<< metal1 >>
rect -196 1281 196 1287
rect -196 1247 -184 1281
rect 184 1247 196 1281
rect -196 1241 196 1247
rect -252 1188 -206 1200
rect -252 -1188 -246 1188
rect -212 -1188 -206 1188
rect -252 -1200 -206 -1188
rect 206 1188 252 1200
rect 206 -1188 212 1188
rect 246 -1188 252 1188
rect 206 -1200 252 -1188
rect -196 -1247 196 -1241
rect -196 -1281 -184 -1247
rect 184 -1281 196 -1247
rect -196 -1287 196 -1281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 12.0 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
