magic
tech sky130A
magscale 1 2
timestamp 1681339707
<< nwell >>
rect -4828 7260 -2290 8460
rect 570 7310 3108 8472
rect 6940 7310 9478 8472
rect 13310 7310 15848 8472
rect 19680 7310 22218 8472
rect 28938 7310 31476 8472
<< pmoslvt >>
rect -4668 7360 -4598 8360
rect -4540 7360 -4470 8360
rect -4264 7360 -4194 8360
rect -4136 7360 -4066 8360
rect -3860 7360 -3790 8360
rect -3732 7360 -3662 8360
rect -3456 7360 -3386 8360
rect -3328 7360 -3258 8360
rect -3052 7360 -2982 8360
rect -2924 7360 -2854 8360
rect -2648 7360 -2578 8360
rect -2520 7360 -2450 8360
rect 730 7410 800 8410
rect 858 7410 928 8410
rect 1134 7410 1204 8410
rect 1262 7410 1332 8410
rect 1538 7410 1608 8410
rect 1666 7410 1736 8410
rect 1942 7410 2012 8410
rect 2070 7410 2140 8410
rect 2346 7410 2416 8410
rect 2474 7410 2544 8410
rect 2750 7410 2820 8410
rect 2878 7410 2948 8410
rect 7100 7410 7170 8410
rect 7228 7410 7298 8410
rect 7504 7410 7574 8410
rect 7632 7410 7702 8410
rect 7908 7410 7978 8410
rect 8036 7410 8106 8410
rect 8312 7410 8382 8410
rect 8440 7410 8510 8410
rect 8716 7410 8786 8410
rect 8844 7410 8914 8410
rect 9120 7410 9190 8410
rect 9248 7410 9318 8410
rect 13470 7410 13540 8410
rect 13598 7410 13668 8410
rect 13874 7410 13944 8410
rect 14002 7410 14072 8410
rect 14278 7410 14348 8410
rect 14406 7410 14476 8410
rect 14682 7410 14752 8410
rect 14810 7410 14880 8410
rect 15086 7410 15156 8410
rect 15214 7410 15284 8410
rect 15490 7410 15560 8410
rect 15618 7410 15688 8410
rect 19840 7410 19910 8410
rect 19968 7410 20038 8410
rect 20244 7410 20314 8410
rect 20372 7410 20442 8410
rect 20648 7410 20718 8410
rect 20776 7410 20846 8410
rect 21052 7410 21122 8410
rect 21180 7410 21250 8410
rect 21456 7410 21526 8410
rect 21584 7410 21654 8410
rect 21860 7410 21930 8410
rect 21988 7410 22058 8410
rect 29098 7410 29168 8410
rect 29226 7410 29296 8410
rect 29502 7410 29572 8410
rect 29630 7410 29700 8410
rect 29906 7410 29976 8410
rect 30034 7410 30104 8410
rect 30310 7410 30380 8410
rect 30438 7410 30508 8410
rect 30714 7410 30784 8410
rect 30842 7410 30912 8410
rect 31118 7410 31188 8410
rect 31246 7410 31316 8410
<< nmoslvt >>
rect -4464 5884 -4428 6884
rect -4370 5884 -4334 6884
rect -4128 5884 -4092 6884
rect -4034 5884 -3998 6884
rect -3792 5884 -3756 6884
rect -3698 5884 -3662 6884
rect -3456 5884 -3420 6884
rect -3362 5884 -3326 6884
rect -3120 5884 -3084 6884
rect -3026 5884 -2990 6884
rect -2784 5884 -2748 6884
rect -2690 5884 -2654 6884
rect 934 5934 970 6934
rect 1028 5934 1064 6934
rect 1270 5934 1306 6934
rect 1364 5934 1400 6934
rect 1606 5934 1642 6934
rect 1700 5934 1736 6934
rect 1942 5934 1978 6934
rect 2036 5934 2072 6934
rect 2278 5934 2314 6934
rect 2372 5934 2408 6934
rect 2614 5934 2650 6934
rect 2708 5934 2744 6934
rect 7304 5934 7340 6934
rect 7398 5934 7434 6934
rect 7640 5934 7676 6934
rect 7734 5934 7770 6934
rect 7976 5934 8012 6934
rect 8070 5934 8106 6934
rect 8312 5934 8348 6934
rect 8406 5934 8442 6934
rect 8648 5934 8684 6934
rect 8742 5934 8778 6934
rect 8984 5934 9020 6934
rect 9078 5934 9114 6934
rect 13674 5934 13710 6934
rect 13768 5934 13804 6934
rect 14010 5934 14046 6934
rect 14104 5934 14140 6934
rect 14346 5934 14382 6934
rect 14440 5934 14476 6934
rect 14682 5934 14718 6934
rect 14776 5934 14812 6934
rect 15018 5934 15054 6934
rect 15112 5934 15148 6934
rect 15354 5934 15390 6934
rect 15448 5934 15484 6934
rect 20044 5934 20080 6934
rect 20138 5934 20174 6934
rect 20380 5934 20416 6934
rect 20474 5934 20510 6934
rect 20716 5934 20752 6934
rect 20810 5934 20846 6934
rect 21052 5934 21088 6934
rect 21146 5934 21182 6934
rect 21388 5934 21424 6934
rect 21482 5934 21518 6934
rect 21724 5934 21760 6934
rect 21818 5934 21854 6934
rect 29302 5934 29338 6934
rect 29396 5934 29432 6934
rect 29638 5934 29674 6934
rect 29732 5934 29768 6934
rect 29974 5934 30010 6934
rect 30068 5934 30104 6934
rect 30310 5934 30346 6934
rect 30404 5934 30440 6934
rect 30646 5934 30682 6934
rect 30740 5934 30776 6934
rect 30982 5934 31018 6934
rect 31076 5934 31112 6934
<< ndiff >>
rect -4524 6872 -4464 6884
rect -4524 5896 -4510 6872
rect -4476 5896 -4464 6872
rect -4524 5884 -4464 5896
rect -4428 6872 -4370 6884
rect -4428 5896 -4416 6872
rect -4382 5896 -4370 6872
rect -4428 5884 -4370 5896
rect -4334 6872 -4274 6884
rect -4334 5896 -4322 6872
rect -4288 5896 -4274 6872
rect -4188 6872 -4128 6884
rect -4334 5884 -4274 5896
rect -4188 5896 -4174 6872
rect -4140 5896 -4128 6872
rect -4188 5884 -4128 5896
rect -4092 6872 -4034 6884
rect -4092 5896 -4080 6872
rect -4046 5896 -4034 6872
rect -4092 5884 -4034 5896
rect -3998 6872 -3938 6884
rect -3998 5896 -3986 6872
rect -3952 5896 -3938 6872
rect -3852 6872 -3792 6884
rect -3998 5884 -3938 5896
rect -3852 5896 -3838 6872
rect -3804 5896 -3792 6872
rect -3852 5884 -3792 5896
rect -3756 6872 -3698 6884
rect -3756 5896 -3744 6872
rect -3710 5896 -3698 6872
rect -3756 5884 -3698 5896
rect -3662 6872 -3602 6884
rect -3662 5896 -3650 6872
rect -3616 5896 -3602 6872
rect -3516 6872 -3456 6884
rect -3662 5884 -3602 5896
rect -3516 5896 -3502 6872
rect -3468 5896 -3456 6872
rect -3516 5884 -3456 5896
rect -3420 6872 -3362 6884
rect -3420 5896 -3408 6872
rect -3374 5896 -3362 6872
rect -3420 5884 -3362 5896
rect -3326 6872 -3266 6884
rect -3326 5896 -3314 6872
rect -3280 5896 -3266 6872
rect -3180 6872 -3120 6884
rect -3326 5884 -3266 5896
rect -3180 5896 -3166 6872
rect -3132 5896 -3120 6872
rect -3180 5884 -3120 5896
rect -3084 6872 -3026 6884
rect -3084 5896 -3072 6872
rect -3038 5896 -3026 6872
rect -3084 5884 -3026 5896
rect -2990 6872 -2930 6884
rect -2990 5896 -2978 6872
rect -2944 5896 -2930 6872
rect -2844 6872 -2784 6884
rect -2990 5884 -2930 5896
rect -2844 5896 -2830 6872
rect -2796 5896 -2784 6872
rect -2844 5884 -2784 5896
rect -2748 6872 -2690 6884
rect -2748 5896 -2736 6872
rect -2702 5896 -2690 6872
rect -2748 5884 -2690 5896
rect -2654 6872 -2594 6884
rect -2654 5896 -2642 6872
rect -2608 5896 -2594 6872
rect -2654 5884 -2594 5896
rect 874 6922 934 6934
rect 874 5946 888 6922
rect 922 5946 934 6922
rect 874 5934 934 5946
rect 970 6922 1028 6934
rect 970 5946 982 6922
rect 1016 5946 1028 6922
rect 970 5934 1028 5946
rect 1064 6922 1124 6934
rect 1064 5946 1076 6922
rect 1110 5946 1124 6922
rect 1210 6922 1270 6934
rect 1064 5934 1124 5946
rect 1210 5946 1224 6922
rect 1258 5946 1270 6922
rect 1210 5934 1270 5946
rect 1306 6922 1364 6934
rect 1306 5946 1318 6922
rect 1352 5946 1364 6922
rect 1306 5934 1364 5946
rect 1400 6922 1460 6934
rect 1400 5946 1412 6922
rect 1446 5946 1460 6922
rect 1546 6922 1606 6934
rect 1400 5934 1460 5946
rect 1546 5946 1560 6922
rect 1594 5946 1606 6922
rect 1546 5934 1606 5946
rect 1642 6922 1700 6934
rect 1642 5946 1654 6922
rect 1688 5946 1700 6922
rect 1642 5934 1700 5946
rect 1736 6922 1796 6934
rect 1736 5946 1748 6922
rect 1782 5946 1796 6922
rect 1882 6922 1942 6934
rect 1736 5934 1796 5946
rect 1882 5946 1896 6922
rect 1930 5946 1942 6922
rect 1882 5934 1942 5946
rect 1978 6922 2036 6934
rect 1978 5946 1990 6922
rect 2024 5946 2036 6922
rect 1978 5934 2036 5946
rect 2072 6922 2132 6934
rect 2072 5946 2084 6922
rect 2118 5946 2132 6922
rect 2218 6922 2278 6934
rect 2072 5934 2132 5946
rect 2218 5946 2232 6922
rect 2266 5946 2278 6922
rect 2218 5934 2278 5946
rect 2314 6922 2372 6934
rect 2314 5946 2326 6922
rect 2360 5946 2372 6922
rect 2314 5934 2372 5946
rect 2408 6922 2468 6934
rect 2408 5946 2420 6922
rect 2454 5946 2468 6922
rect 2554 6922 2614 6934
rect 2408 5934 2468 5946
rect 2554 5946 2568 6922
rect 2602 5946 2614 6922
rect 2554 5934 2614 5946
rect 2650 6922 2708 6934
rect 2650 5946 2662 6922
rect 2696 5946 2708 6922
rect 2650 5934 2708 5946
rect 2744 6922 2804 6934
rect 2744 5946 2756 6922
rect 2790 5946 2804 6922
rect 2744 5934 2804 5946
rect 7244 6922 7304 6934
rect 7244 5946 7258 6922
rect 7292 5946 7304 6922
rect 7244 5934 7304 5946
rect 7340 6922 7398 6934
rect 7340 5946 7352 6922
rect 7386 5946 7398 6922
rect 7340 5934 7398 5946
rect 7434 6922 7494 6934
rect 7434 5946 7446 6922
rect 7480 5946 7494 6922
rect 7580 6922 7640 6934
rect 7434 5934 7494 5946
rect 7580 5946 7594 6922
rect 7628 5946 7640 6922
rect 7580 5934 7640 5946
rect 7676 6922 7734 6934
rect 7676 5946 7688 6922
rect 7722 5946 7734 6922
rect 7676 5934 7734 5946
rect 7770 6922 7830 6934
rect 7770 5946 7782 6922
rect 7816 5946 7830 6922
rect 7916 6922 7976 6934
rect 7770 5934 7830 5946
rect 7916 5946 7930 6922
rect 7964 5946 7976 6922
rect 7916 5934 7976 5946
rect 8012 6922 8070 6934
rect 8012 5946 8024 6922
rect 8058 5946 8070 6922
rect 8012 5934 8070 5946
rect 8106 6922 8166 6934
rect 8106 5946 8118 6922
rect 8152 5946 8166 6922
rect 8252 6922 8312 6934
rect 8106 5934 8166 5946
rect 8252 5946 8266 6922
rect 8300 5946 8312 6922
rect 8252 5934 8312 5946
rect 8348 6922 8406 6934
rect 8348 5946 8360 6922
rect 8394 5946 8406 6922
rect 8348 5934 8406 5946
rect 8442 6922 8502 6934
rect 8442 5946 8454 6922
rect 8488 5946 8502 6922
rect 8588 6922 8648 6934
rect 8442 5934 8502 5946
rect 8588 5946 8602 6922
rect 8636 5946 8648 6922
rect 8588 5934 8648 5946
rect 8684 6922 8742 6934
rect 8684 5946 8696 6922
rect 8730 5946 8742 6922
rect 8684 5934 8742 5946
rect 8778 6922 8838 6934
rect 8778 5946 8790 6922
rect 8824 5946 8838 6922
rect 8924 6922 8984 6934
rect 8778 5934 8838 5946
rect 8924 5946 8938 6922
rect 8972 5946 8984 6922
rect 8924 5934 8984 5946
rect 9020 6922 9078 6934
rect 9020 5946 9032 6922
rect 9066 5946 9078 6922
rect 9020 5934 9078 5946
rect 9114 6922 9174 6934
rect 9114 5946 9126 6922
rect 9160 5946 9174 6922
rect 9114 5934 9174 5946
rect 13614 6922 13674 6934
rect 13614 5946 13628 6922
rect 13662 5946 13674 6922
rect 13614 5934 13674 5946
rect 13710 6922 13768 6934
rect 13710 5946 13722 6922
rect 13756 5946 13768 6922
rect 13710 5934 13768 5946
rect 13804 6922 13864 6934
rect 13804 5946 13816 6922
rect 13850 5946 13864 6922
rect 13950 6922 14010 6934
rect 13804 5934 13864 5946
rect 13950 5946 13964 6922
rect 13998 5946 14010 6922
rect 13950 5934 14010 5946
rect 14046 6922 14104 6934
rect 14046 5946 14058 6922
rect 14092 5946 14104 6922
rect 14046 5934 14104 5946
rect 14140 6922 14200 6934
rect 14140 5946 14152 6922
rect 14186 5946 14200 6922
rect 14286 6922 14346 6934
rect 14140 5934 14200 5946
rect 14286 5946 14300 6922
rect 14334 5946 14346 6922
rect 14286 5934 14346 5946
rect 14382 6922 14440 6934
rect 14382 5946 14394 6922
rect 14428 5946 14440 6922
rect 14382 5934 14440 5946
rect 14476 6922 14536 6934
rect 14476 5946 14488 6922
rect 14522 5946 14536 6922
rect 14622 6922 14682 6934
rect 14476 5934 14536 5946
rect 14622 5946 14636 6922
rect 14670 5946 14682 6922
rect 14622 5934 14682 5946
rect 14718 6922 14776 6934
rect 14718 5946 14730 6922
rect 14764 5946 14776 6922
rect 14718 5934 14776 5946
rect 14812 6922 14872 6934
rect 14812 5946 14824 6922
rect 14858 5946 14872 6922
rect 14958 6922 15018 6934
rect 14812 5934 14872 5946
rect 14958 5946 14972 6922
rect 15006 5946 15018 6922
rect 14958 5934 15018 5946
rect 15054 6922 15112 6934
rect 15054 5946 15066 6922
rect 15100 5946 15112 6922
rect 15054 5934 15112 5946
rect 15148 6922 15208 6934
rect 15148 5946 15160 6922
rect 15194 5946 15208 6922
rect 15294 6922 15354 6934
rect 15148 5934 15208 5946
rect 15294 5946 15308 6922
rect 15342 5946 15354 6922
rect 15294 5934 15354 5946
rect 15390 6922 15448 6934
rect 15390 5946 15402 6922
rect 15436 5946 15448 6922
rect 15390 5934 15448 5946
rect 15484 6922 15544 6934
rect 15484 5946 15496 6922
rect 15530 5946 15544 6922
rect 15484 5934 15544 5946
rect 19984 6922 20044 6934
rect 19984 5946 19998 6922
rect 20032 5946 20044 6922
rect 19984 5934 20044 5946
rect 20080 6922 20138 6934
rect 20080 5946 20092 6922
rect 20126 5946 20138 6922
rect 20080 5934 20138 5946
rect 20174 6922 20234 6934
rect 20174 5946 20186 6922
rect 20220 5946 20234 6922
rect 20320 6922 20380 6934
rect 20174 5934 20234 5946
rect 20320 5946 20334 6922
rect 20368 5946 20380 6922
rect 20320 5934 20380 5946
rect 20416 6922 20474 6934
rect 20416 5946 20428 6922
rect 20462 5946 20474 6922
rect 20416 5934 20474 5946
rect 20510 6922 20570 6934
rect 20510 5946 20522 6922
rect 20556 5946 20570 6922
rect 20656 6922 20716 6934
rect 20510 5934 20570 5946
rect 20656 5946 20670 6922
rect 20704 5946 20716 6922
rect 20656 5934 20716 5946
rect 20752 6922 20810 6934
rect 20752 5946 20764 6922
rect 20798 5946 20810 6922
rect 20752 5934 20810 5946
rect 20846 6922 20906 6934
rect 20846 5946 20858 6922
rect 20892 5946 20906 6922
rect 20992 6922 21052 6934
rect 20846 5934 20906 5946
rect 20992 5946 21006 6922
rect 21040 5946 21052 6922
rect 20992 5934 21052 5946
rect 21088 6922 21146 6934
rect 21088 5946 21100 6922
rect 21134 5946 21146 6922
rect 21088 5934 21146 5946
rect 21182 6922 21242 6934
rect 21182 5946 21194 6922
rect 21228 5946 21242 6922
rect 21328 6922 21388 6934
rect 21182 5934 21242 5946
rect 21328 5946 21342 6922
rect 21376 5946 21388 6922
rect 21328 5934 21388 5946
rect 21424 6922 21482 6934
rect 21424 5946 21436 6922
rect 21470 5946 21482 6922
rect 21424 5934 21482 5946
rect 21518 6922 21578 6934
rect 21518 5946 21530 6922
rect 21564 5946 21578 6922
rect 21664 6922 21724 6934
rect 21518 5934 21578 5946
rect 21664 5946 21678 6922
rect 21712 5946 21724 6922
rect 21664 5934 21724 5946
rect 21760 6922 21818 6934
rect 21760 5946 21772 6922
rect 21806 5946 21818 6922
rect 21760 5934 21818 5946
rect 21854 6922 21914 6934
rect 21854 5946 21866 6922
rect 21900 5946 21914 6922
rect 21854 5934 21914 5946
rect 29242 6922 29302 6934
rect 29242 5946 29256 6922
rect 29290 5946 29302 6922
rect 29242 5934 29302 5946
rect 29338 6922 29396 6934
rect 29338 5946 29350 6922
rect 29384 5946 29396 6922
rect 29338 5934 29396 5946
rect 29432 6922 29492 6934
rect 29432 5946 29444 6922
rect 29478 5946 29492 6922
rect 29578 6922 29638 6934
rect 29432 5934 29492 5946
rect 29578 5946 29592 6922
rect 29626 5946 29638 6922
rect 29578 5934 29638 5946
rect 29674 6922 29732 6934
rect 29674 5946 29686 6922
rect 29720 5946 29732 6922
rect 29674 5934 29732 5946
rect 29768 6922 29828 6934
rect 29768 5946 29780 6922
rect 29814 5946 29828 6922
rect 29914 6922 29974 6934
rect 29768 5934 29828 5946
rect 29914 5946 29928 6922
rect 29962 5946 29974 6922
rect 29914 5934 29974 5946
rect 30010 6922 30068 6934
rect 30010 5946 30022 6922
rect 30056 5946 30068 6922
rect 30010 5934 30068 5946
rect 30104 6922 30164 6934
rect 30104 5946 30116 6922
rect 30150 5946 30164 6922
rect 30250 6922 30310 6934
rect 30104 5934 30164 5946
rect 30250 5946 30264 6922
rect 30298 5946 30310 6922
rect 30250 5934 30310 5946
rect 30346 6922 30404 6934
rect 30346 5946 30358 6922
rect 30392 5946 30404 6922
rect 30346 5934 30404 5946
rect 30440 6922 30500 6934
rect 30440 5946 30452 6922
rect 30486 5946 30500 6922
rect 30586 6922 30646 6934
rect 30440 5934 30500 5946
rect 30586 5946 30600 6922
rect 30634 5946 30646 6922
rect 30586 5934 30646 5946
rect 30682 6922 30740 6934
rect 30682 5946 30694 6922
rect 30728 5946 30740 6922
rect 30682 5934 30740 5946
rect 30776 6922 30836 6934
rect 30776 5946 30788 6922
rect 30822 5946 30836 6922
rect 30922 6922 30982 6934
rect 30776 5934 30836 5946
rect 30922 5946 30936 6922
rect 30970 5946 30982 6922
rect 30922 5934 30982 5946
rect 31018 6922 31076 6934
rect 31018 5946 31030 6922
rect 31064 5946 31076 6922
rect 31018 5934 31076 5946
rect 31112 6922 31172 6934
rect 31112 5946 31124 6922
rect 31158 5946 31172 6922
rect 31112 5934 31172 5946
<< pdiff >>
rect -4728 8348 -4668 8360
rect -4728 7372 -4714 8348
rect -4680 7372 -4668 8348
rect -4728 7360 -4668 7372
rect -4598 8348 -4540 8360
rect -4598 7372 -4586 8348
rect -4552 7372 -4540 8348
rect -4598 7360 -4540 7372
rect -4470 8348 -4410 8360
rect -4470 7372 -4458 8348
rect -4424 7372 -4410 8348
rect -4324 8348 -4264 8360
rect -4470 7360 -4410 7372
rect -4324 7372 -4310 8348
rect -4276 7372 -4264 8348
rect -4324 7360 -4264 7372
rect -4194 8348 -4136 8360
rect -4194 7372 -4182 8348
rect -4148 7372 -4136 8348
rect -4194 7360 -4136 7372
rect -4066 8348 -4006 8360
rect -4066 7372 -4054 8348
rect -4020 7372 -4006 8348
rect -3920 8348 -3860 8360
rect -4066 7360 -4006 7372
rect -3920 7372 -3906 8348
rect -3872 7372 -3860 8348
rect -3920 7360 -3860 7372
rect -3790 8348 -3732 8360
rect -3790 7372 -3778 8348
rect -3744 7372 -3732 8348
rect -3790 7360 -3732 7372
rect -3662 8348 -3602 8360
rect -3662 7372 -3650 8348
rect -3616 7372 -3602 8348
rect -3516 8348 -3456 8360
rect -3662 7360 -3602 7372
rect -3516 7372 -3502 8348
rect -3468 7372 -3456 8348
rect -3516 7360 -3456 7372
rect -3386 8348 -3328 8360
rect -3386 7372 -3374 8348
rect -3340 7372 -3328 8348
rect -3386 7360 -3328 7372
rect -3258 8348 -3198 8360
rect -3258 7372 -3246 8348
rect -3212 7372 -3198 8348
rect -3112 8348 -3052 8360
rect -3258 7360 -3198 7372
rect -3112 7372 -3098 8348
rect -3064 7372 -3052 8348
rect -3112 7360 -3052 7372
rect -2982 8348 -2924 8360
rect -2982 7372 -2970 8348
rect -2936 7372 -2924 8348
rect -2982 7360 -2924 7372
rect -2854 8348 -2794 8360
rect -2854 7372 -2842 8348
rect -2808 7372 -2794 8348
rect -2708 8348 -2648 8360
rect -2854 7360 -2794 7372
rect -2708 7372 -2694 8348
rect -2660 7372 -2648 8348
rect -2708 7360 -2648 7372
rect -2578 8348 -2520 8360
rect -2578 7372 -2566 8348
rect -2532 7372 -2520 8348
rect -2578 7360 -2520 7372
rect -2450 8348 -2390 8360
rect -2450 7372 -2438 8348
rect -2404 7372 -2390 8348
rect -2450 7360 -2390 7372
rect 670 8398 730 8410
rect 670 7422 684 8398
rect 718 7422 730 8398
rect 670 7410 730 7422
rect 800 8398 858 8410
rect 800 7422 812 8398
rect 846 7422 858 8398
rect 800 7410 858 7422
rect 928 8398 988 8410
rect 928 7422 940 8398
rect 974 7422 988 8398
rect 1074 8398 1134 8410
rect 928 7410 988 7422
rect 1074 7422 1088 8398
rect 1122 7422 1134 8398
rect 1074 7410 1134 7422
rect 1204 8398 1262 8410
rect 1204 7422 1216 8398
rect 1250 7422 1262 8398
rect 1204 7410 1262 7422
rect 1332 8398 1392 8410
rect 1332 7422 1344 8398
rect 1378 7422 1392 8398
rect 1478 8398 1538 8410
rect 1332 7410 1392 7422
rect 1478 7422 1492 8398
rect 1526 7422 1538 8398
rect 1478 7410 1538 7422
rect 1608 8398 1666 8410
rect 1608 7422 1620 8398
rect 1654 7422 1666 8398
rect 1608 7410 1666 7422
rect 1736 8398 1796 8410
rect 1736 7422 1748 8398
rect 1782 7422 1796 8398
rect 1882 8398 1942 8410
rect 1736 7410 1796 7422
rect 1882 7422 1896 8398
rect 1930 7422 1942 8398
rect 1882 7410 1942 7422
rect 2012 8398 2070 8410
rect 2012 7422 2024 8398
rect 2058 7422 2070 8398
rect 2012 7410 2070 7422
rect 2140 8398 2200 8410
rect 2140 7422 2152 8398
rect 2186 7422 2200 8398
rect 2286 8398 2346 8410
rect 2140 7410 2200 7422
rect 2286 7422 2300 8398
rect 2334 7422 2346 8398
rect 2286 7410 2346 7422
rect 2416 8398 2474 8410
rect 2416 7422 2428 8398
rect 2462 7422 2474 8398
rect 2416 7410 2474 7422
rect 2544 8398 2604 8410
rect 2544 7422 2556 8398
rect 2590 7422 2604 8398
rect 2690 8398 2750 8410
rect 2544 7410 2604 7422
rect 2690 7422 2704 8398
rect 2738 7422 2750 8398
rect 2690 7410 2750 7422
rect 2820 8398 2878 8410
rect 2820 7422 2832 8398
rect 2866 7422 2878 8398
rect 2820 7410 2878 7422
rect 2948 8398 3008 8410
rect 2948 7422 2960 8398
rect 2994 7422 3008 8398
rect 2948 7410 3008 7422
rect 7040 8398 7100 8410
rect 7040 7422 7054 8398
rect 7088 7422 7100 8398
rect 7040 7410 7100 7422
rect 7170 8398 7228 8410
rect 7170 7422 7182 8398
rect 7216 7422 7228 8398
rect 7170 7410 7228 7422
rect 7298 8398 7358 8410
rect 7298 7422 7310 8398
rect 7344 7422 7358 8398
rect 7444 8398 7504 8410
rect 7298 7410 7358 7422
rect 7444 7422 7458 8398
rect 7492 7422 7504 8398
rect 7444 7410 7504 7422
rect 7574 8398 7632 8410
rect 7574 7422 7586 8398
rect 7620 7422 7632 8398
rect 7574 7410 7632 7422
rect 7702 8398 7762 8410
rect 7702 7422 7714 8398
rect 7748 7422 7762 8398
rect 7848 8398 7908 8410
rect 7702 7410 7762 7422
rect 7848 7422 7862 8398
rect 7896 7422 7908 8398
rect 7848 7410 7908 7422
rect 7978 8398 8036 8410
rect 7978 7422 7990 8398
rect 8024 7422 8036 8398
rect 7978 7410 8036 7422
rect 8106 8398 8166 8410
rect 8106 7422 8118 8398
rect 8152 7422 8166 8398
rect 8252 8398 8312 8410
rect 8106 7410 8166 7422
rect 8252 7422 8266 8398
rect 8300 7422 8312 8398
rect 8252 7410 8312 7422
rect 8382 8398 8440 8410
rect 8382 7422 8394 8398
rect 8428 7422 8440 8398
rect 8382 7410 8440 7422
rect 8510 8398 8570 8410
rect 8510 7422 8522 8398
rect 8556 7422 8570 8398
rect 8656 8398 8716 8410
rect 8510 7410 8570 7422
rect 8656 7422 8670 8398
rect 8704 7422 8716 8398
rect 8656 7410 8716 7422
rect 8786 8398 8844 8410
rect 8786 7422 8798 8398
rect 8832 7422 8844 8398
rect 8786 7410 8844 7422
rect 8914 8398 8974 8410
rect 8914 7422 8926 8398
rect 8960 7422 8974 8398
rect 9060 8398 9120 8410
rect 8914 7410 8974 7422
rect 9060 7422 9074 8398
rect 9108 7422 9120 8398
rect 9060 7410 9120 7422
rect 9190 8398 9248 8410
rect 9190 7422 9202 8398
rect 9236 7422 9248 8398
rect 9190 7410 9248 7422
rect 9318 8398 9378 8410
rect 9318 7422 9330 8398
rect 9364 7422 9378 8398
rect 9318 7410 9378 7422
rect 13410 8398 13470 8410
rect 13410 7422 13424 8398
rect 13458 7422 13470 8398
rect 13410 7410 13470 7422
rect 13540 8398 13598 8410
rect 13540 7422 13552 8398
rect 13586 7422 13598 8398
rect 13540 7410 13598 7422
rect 13668 8398 13728 8410
rect 13668 7422 13680 8398
rect 13714 7422 13728 8398
rect 13814 8398 13874 8410
rect 13668 7410 13728 7422
rect 13814 7422 13828 8398
rect 13862 7422 13874 8398
rect 13814 7410 13874 7422
rect 13944 8398 14002 8410
rect 13944 7422 13956 8398
rect 13990 7422 14002 8398
rect 13944 7410 14002 7422
rect 14072 8398 14132 8410
rect 14072 7422 14084 8398
rect 14118 7422 14132 8398
rect 14218 8398 14278 8410
rect 14072 7410 14132 7422
rect 14218 7422 14232 8398
rect 14266 7422 14278 8398
rect 14218 7410 14278 7422
rect 14348 8398 14406 8410
rect 14348 7422 14360 8398
rect 14394 7422 14406 8398
rect 14348 7410 14406 7422
rect 14476 8398 14536 8410
rect 14476 7422 14488 8398
rect 14522 7422 14536 8398
rect 14622 8398 14682 8410
rect 14476 7410 14536 7422
rect 14622 7422 14636 8398
rect 14670 7422 14682 8398
rect 14622 7410 14682 7422
rect 14752 8398 14810 8410
rect 14752 7422 14764 8398
rect 14798 7422 14810 8398
rect 14752 7410 14810 7422
rect 14880 8398 14940 8410
rect 14880 7422 14892 8398
rect 14926 7422 14940 8398
rect 15026 8398 15086 8410
rect 14880 7410 14940 7422
rect 15026 7422 15040 8398
rect 15074 7422 15086 8398
rect 15026 7410 15086 7422
rect 15156 8398 15214 8410
rect 15156 7422 15168 8398
rect 15202 7422 15214 8398
rect 15156 7410 15214 7422
rect 15284 8398 15344 8410
rect 15284 7422 15296 8398
rect 15330 7422 15344 8398
rect 15430 8398 15490 8410
rect 15284 7410 15344 7422
rect 15430 7422 15444 8398
rect 15478 7422 15490 8398
rect 15430 7410 15490 7422
rect 15560 8398 15618 8410
rect 15560 7422 15572 8398
rect 15606 7422 15618 8398
rect 15560 7410 15618 7422
rect 15688 8398 15748 8410
rect 15688 7422 15700 8398
rect 15734 7422 15748 8398
rect 15688 7410 15748 7422
rect 19780 8398 19840 8410
rect 19780 7422 19794 8398
rect 19828 7422 19840 8398
rect 19780 7410 19840 7422
rect 19910 8398 19968 8410
rect 19910 7422 19922 8398
rect 19956 7422 19968 8398
rect 19910 7410 19968 7422
rect 20038 8398 20098 8410
rect 20038 7422 20050 8398
rect 20084 7422 20098 8398
rect 20184 8398 20244 8410
rect 20038 7410 20098 7422
rect 20184 7422 20198 8398
rect 20232 7422 20244 8398
rect 20184 7410 20244 7422
rect 20314 8398 20372 8410
rect 20314 7422 20326 8398
rect 20360 7422 20372 8398
rect 20314 7410 20372 7422
rect 20442 8398 20502 8410
rect 20442 7422 20454 8398
rect 20488 7422 20502 8398
rect 20588 8398 20648 8410
rect 20442 7410 20502 7422
rect 20588 7422 20602 8398
rect 20636 7422 20648 8398
rect 20588 7410 20648 7422
rect 20718 8398 20776 8410
rect 20718 7422 20730 8398
rect 20764 7422 20776 8398
rect 20718 7410 20776 7422
rect 20846 8398 20906 8410
rect 20846 7422 20858 8398
rect 20892 7422 20906 8398
rect 20992 8398 21052 8410
rect 20846 7410 20906 7422
rect 20992 7422 21006 8398
rect 21040 7422 21052 8398
rect 20992 7410 21052 7422
rect 21122 8398 21180 8410
rect 21122 7422 21134 8398
rect 21168 7422 21180 8398
rect 21122 7410 21180 7422
rect 21250 8398 21310 8410
rect 21250 7422 21262 8398
rect 21296 7422 21310 8398
rect 21396 8398 21456 8410
rect 21250 7410 21310 7422
rect 21396 7422 21410 8398
rect 21444 7422 21456 8398
rect 21396 7410 21456 7422
rect 21526 8398 21584 8410
rect 21526 7422 21538 8398
rect 21572 7422 21584 8398
rect 21526 7410 21584 7422
rect 21654 8398 21714 8410
rect 21654 7422 21666 8398
rect 21700 7422 21714 8398
rect 21800 8398 21860 8410
rect 21654 7410 21714 7422
rect 21800 7422 21814 8398
rect 21848 7422 21860 8398
rect 21800 7410 21860 7422
rect 21930 8398 21988 8410
rect 21930 7422 21942 8398
rect 21976 7422 21988 8398
rect 21930 7410 21988 7422
rect 22058 8398 22118 8410
rect 22058 7422 22070 8398
rect 22104 7422 22118 8398
rect 22058 7410 22118 7422
rect 29038 8398 29098 8410
rect 29038 7422 29052 8398
rect 29086 7422 29098 8398
rect 29038 7410 29098 7422
rect 29168 8398 29226 8410
rect 29168 7422 29180 8398
rect 29214 7422 29226 8398
rect 29168 7410 29226 7422
rect 29296 8398 29356 8410
rect 29296 7422 29308 8398
rect 29342 7422 29356 8398
rect 29442 8398 29502 8410
rect 29296 7410 29356 7422
rect 29442 7422 29456 8398
rect 29490 7422 29502 8398
rect 29442 7410 29502 7422
rect 29572 8398 29630 8410
rect 29572 7422 29584 8398
rect 29618 7422 29630 8398
rect 29572 7410 29630 7422
rect 29700 8398 29760 8410
rect 29700 7422 29712 8398
rect 29746 7422 29760 8398
rect 29846 8398 29906 8410
rect 29700 7410 29760 7422
rect 29846 7422 29860 8398
rect 29894 7422 29906 8398
rect 29846 7410 29906 7422
rect 29976 8398 30034 8410
rect 29976 7422 29988 8398
rect 30022 7422 30034 8398
rect 29976 7410 30034 7422
rect 30104 8398 30164 8410
rect 30104 7422 30116 8398
rect 30150 7422 30164 8398
rect 30250 8398 30310 8410
rect 30104 7410 30164 7422
rect 30250 7422 30264 8398
rect 30298 7422 30310 8398
rect 30250 7410 30310 7422
rect 30380 8398 30438 8410
rect 30380 7422 30392 8398
rect 30426 7422 30438 8398
rect 30380 7410 30438 7422
rect 30508 8398 30568 8410
rect 30508 7422 30520 8398
rect 30554 7422 30568 8398
rect 30654 8398 30714 8410
rect 30508 7410 30568 7422
rect 30654 7422 30668 8398
rect 30702 7422 30714 8398
rect 30654 7410 30714 7422
rect 30784 8398 30842 8410
rect 30784 7422 30796 8398
rect 30830 7422 30842 8398
rect 30784 7410 30842 7422
rect 30912 8398 30972 8410
rect 30912 7422 30924 8398
rect 30958 7422 30972 8398
rect 31058 8398 31118 8410
rect 30912 7410 30972 7422
rect 31058 7422 31072 8398
rect 31106 7422 31118 8398
rect 31058 7410 31118 7422
rect 31188 8398 31246 8410
rect 31188 7422 31200 8398
rect 31234 7422 31246 8398
rect 31188 7410 31246 7422
rect 31316 8398 31376 8410
rect 31316 7422 31328 8398
rect 31362 7422 31376 8398
rect 31316 7410 31376 7422
<< ndiffc >>
rect -4510 5896 -4476 6872
rect -4416 5896 -4382 6872
rect -4322 5896 -4288 6872
rect -4174 5896 -4140 6872
rect -4080 5896 -4046 6872
rect -3986 5896 -3952 6872
rect -3838 5896 -3804 6872
rect -3744 5896 -3710 6872
rect -3650 5896 -3616 6872
rect -3502 5896 -3468 6872
rect -3408 5896 -3374 6872
rect -3314 5896 -3280 6872
rect -3166 5896 -3132 6872
rect -3072 5896 -3038 6872
rect -2978 5896 -2944 6872
rect -2830 5896 -2796 6872
rect -2736 5896 -2702 6872
rect -2642 5896 -2608 6872
rect 888 5946 922 6922
rect 982 5946 1016 6922
rect 1076 5946 1110 6922
rect 1224 5946 1258 6922
rect 1318 5946 1352 6922
rect 1412 5946 1446 6922
rect 1560 5946 1594 6922
rect 1654 5946 1688 6922
rect 1748 5946 1782 6922
rect 1896 5946 1930 6922
rect 1990 5946 2024 6922
rect 2084 5946 2118 6922
rect 2232 5946 2266 6922
rect 2326 5946 2360 6922
rect 2420 5946 2454 6922
rect 2568 5946 2602 6922
rect 2662 5946 2696 6922
rect 2756 5946 2790 6922
rect 7258 5946 7292 6922
rect 7352 5946 7386 6922
rect 7446 5946 7480 6922
rect 7594 5946 7628 6922
rect 7688 5946 7722 6922
rect 7782 5946 7816 6922
rect 7930 5946 7964 6922
rect 8024 5946 8058 6922
rect 8118 5946 8152 6922
rect 8266 5946 8300 6922
rect 8360 5946 8394 6922
rect 8454 5946 8488 6922
rect 8602 5946 8636 6922
rect 8696 5946 8730 6922
rect 8790 5946 8824 6922
rect 8938 5946 8972 6922
rect 9032 5946 9066 6922
rect 9126 5946 9160 6922
rect 13628 5946 13662 6922
rect 13722 5946 13756 6922
rect 13816 5946 13850 6922
rect 13964 5946 13998 6922
rect 14058 5946 14092 6922
rect 14152 5946 14186 6922
rect 14300 5946 14334 6922
rect 14394 5946 14428 6922
rect 14488 5946 14522 6922
rect 14636 5946 14670 6922
rect 14730 5946 14764 6922
rect 14824 5946 14858 6922
rect 14972 5946 15006 6922
rect 15066 5946 15100 6922
rect 15160 5946 15194 6922
rect 15308 5946 15342 6922
rect 15402 5946 15436 6922
rect 15496 5946 15530 6922
rect 19998 5946 20032 6922
rect 20092 5946 20126 6922
rect 20186 5946 20220 6922
rect 20334 5946 20368 6922
rect 20428 5946 20462 6922
rect 20522 5946 20556 6922
rect 20670 5946 20704 6922
rect 20764 5946 20798 6922
rect 20858 5946 20892 6922
rect 21006 5946 21040 6922
rect 21100 5946 21134 6922
rect 21194 5946 21228 6922
rect 21342 5946 21376 6922
rect 21436 5946 21470 6922
rect 21530 5946 21564 6922
rect 21678 5946 21712 6922
rect 21772 5946 21806 6922
rect 21866 5946 21900 6922
rect 29256 5946 29290 6922
rect 29350 5946 29384 6922
rect 29444 5946 29478 6922
rect 29592 5946 29626 6922
rect 29686 5946 29720 6922
rect 29780 5946 29814 6922
rect 29928 5946 29962 6922
rect 30022 5946 30056 6922
rect 30116 5946 30150 6922
rect 30264 5946 30298 6922
rect 30358 5946 30392 6922
rect 30452 5946 30486 6922
rect 30600 5946 30634 6922
rect 30694 5946 30728 6922
rect 30788 5946 30822 6922
rect 30936 5946 30970 6922
rect 31030 5946 31064 6922
rect 31124 5946 31158 6922
<< pdiffc >>
rect -4714 7372 -4680 8348
rect -4586 7372 -4552 8348
rect -4458 7372 -4424 8348
rect -4310 7372 -4276 8348
rect -4182 7372 -4148 8348
rect -4054 7372 -4020 8348
rect -3906 7372 -3872 8348
rect -3778 7372 -3744 8348
rect -3650 7372 -3616 8348
rect -3502 7372 -3468 8348
rect -3374 7372 -3340 8348
rect -3246 7372 -3212 8348
rect -3098 7372 -3064 8348
rect -2970 7372 -2936 8348
rect -2842 7372 -2808 8348
rect -2694 7372 -2660 8348
rect -2566 7372 -2532 8348
rect -2438 7372 -2404 8348
rect 684 7422 718 8398
rect 812 7422 846 8398
rect 940 7422 974 8398
rect 1088 7422 1122 8398
rect 1216 7422 1250 8398
rect 1344 7422 1378 8398
rect 1492 7422 1526 8398
rect 1620 7422 1654 8398
rect 1748 7422 1782 8398
rect 1896 7422 1930 8398
rect 2024 7422 2058 8398
rect 2152 7422 2186 8398
rect 2300 7422 2334 8398
rect 2428 7422 2462 8398
rect 2556 7422 2590 8398
rect 2704 7422 2738 8398
rect 2832 7422 2866 8398
rect 2960 7422 2994 8398
rect 7054 7422 7088 8398
rect 7182 7422 7216 8398
rect 7310 7422 7344 8398
rect 7458 7422 7492 8398
rect 7586 7422 7620 8398
rect 7714 7422 7748 8398
rect 7862 7422 7896 8398
rect 7990 7422 8024 8398
rect 8118 7422 8152 8398
rect 8266 7422 8300 8398
rect 8394 7422 8428 8398
rect 8522 7422 8556 8398
rect 8670 7422 8704 8398
rect 8798 7422 8832 8398
rect 8926 7422 8960 8398
rect 9074 7422 9108 8398
rect 9202 7422 9236 8398
rect 9330 7422 9364 8398
rect 13424 7422 13458 8398
rect 13552 7422 13586 8398
rect 13680 7422 13714 8398
rect 13828 7422 13862 8398
rect 13956 7422 13990 8398
rect 14084 7422 14118 8398
rect 14232 7422 14266 8398
rect 14360 7422 14394 8398
rect 14488 7422 14522 8398
rect 14636 7422 14670 8398
rect 14764 7422 14798 8398
rect 14892 7422 14926 8398
rect 15040 7422 15074 8398
rect 15168 7422 15202 8398
rect 15296 7422 15330 8398
rect 15444 7422 15478 8398
rect 15572 7422 15606 8398
rect 15700 7422 15734 8398
rect 19794 7422 19828 8398
rect 19922 7422 19956 8398
rect 20050 7422 20084 8398
rect 20198 7422 20232 8398
rect 20326 7422 20360 8398
rect 20454 7422 20488 8398
rect 20602 7422 20636 8398
rect 20730 7422 20764 8398
rect 20858 7422 20892 8398
rect 21006 7422 21040 8398
rect 21134 7422 21168 8398
rect 21262 7422 21296 8398
rect 21410 7422 21444 8398
rect 21538 7422 21572 8398
rect 21666 7422 21700 8398
rect 21814 7422 21848 8398
rect 21942 7422 21976 8398
rect 22070 7422 22104 8398
rect 29052 7422 29086 8398
rect 29180 7422 29214 8398
rect 29308 7422 29342 8398
rect 29456 7422 29490 8398
rect 29584 7422 29618 8398
rect 29712 7422 29746 8398
rect 29860 7422 29894 8398
rect 29988 7422 30022 8398
rect 30116 7422 30150 8398
rect 30264 7422 30298 8398
rect 30392 7422 30426 8398
rect 30520 7422 30554 8398
rect 30668 7422 30702 8398
rect 30796 7422 30830 8398
rect 30924 7422 30958 8398
rect 31072 7422 31106 8398
rect 31200 7422 31234 8398
rect 31328 7422 31362 8398
<< psubdiff >>
rect -4588 6830 -4524 6884
rect -4588 6796 -4584 6830
rect -4550 6796 -4524 6830
rect -4588 6762 -4524 6796
rect -4588 6728 -4584 6762
rect -4550 6728 -4524 6762
rect -4588 6694 -4524 6728
rect -4588 6660 -4584 6694
rect -4550 6660 -4524 6694
rect -4588 6626 -4524 6660
rect -4588 6592 -4584 6626
rect -4550 6592 -4524 6626
rect -4588 6558 -4524 6592
rect -4588 6524 -4584 6558
rect -4550 6524 -4524 6558
rect -4588 6490 -4524 6524
rect -4588 6456 -4584 6490
rect -4550 6456 -4524 6490
rect -4588 6422 -4524 6456
rect -4588 6388 -4584 6422
rect -4550 6388 -4524 6422
rect -4588 6354 -4524 6388
rect -4588 6320 -4584 6354
rect -4550 6320 -4524 6354
rect -4588 6286 -4524 6320
rect -4588 6252 -4584 6286
rect -4550 6252 -4524 6286
rect -4588 6218 -4524 6252
rect -4588 6184 -4584 6218
rect -4550 6184 -4524 6218
rect -4588 6150 -4524 6184
rect -4588 6116 -4584 6150
rect -4550 6116 -4524 6150
rect -4588 6082 -4524 6116
rect -4588 6048 -4584 6082
rect -4550 6048 -4524 6082
rect -4588 6014 -4524 6048
rect -4588 5980 -4584 6014
rect -4550 5980 -4524 6014
rect -4588 5946 -4524 5980
rect -4588 5912 -4584 5946
rect -4550 5912 -4524 5946
rect -4588 5884 -4524 5912
rect -4274 6856 -4188 6884
rect -4274 6822 -4248 6856
rect -4214 6822 -4188 6856
rect -4274 6788 -4188 6822
rect -4274 6754 -4248 6788
rect -4214 6754 -4188 6788
rect -4274 6720 -4188 6754
rect -4274 6686 -4248 6720
rect -4214 6686 -4188 6720
rect -4274 6652 -4188 6686
rect -4274 6618 -4248 6652
rect -4214 6618 -4188 6652
rect -4274 6584 -4188 6618
rect -4274 6550 -4248 6584
rect -4214 6550 -4188 6584
rect -4274 6516 -4188 6550
rect -4274 6482 -4248 6516
rect -4214 6482 -4188 6516
rect -4274 6448 -4188 6482
rect -4274 6414 -4248 6448
rect -4214 6414 -4188 6448
rect -4274 6380 -4188 6414
rect -4274 6346 -4248 6380
rect -4214 6346 -4188 6380
rect -4274 6312 -4188 6346
rect -4274 6278 -4248 6312
rect -4214 6278 -4188 6312
rect -4274 6244 -4188 6278
rect -4274 6210 -4248 6244
rect -4214 6210 -4188 6244
rect -4274 6176 -4188 6210
rect -4274 6142 -4248 6176
rect -4214 6142 -4188 6176
rect -4274 6108 -4188 6142
rect -4274 6074 -4248 6108
rect -4214 6074 -4188 6108
rect -4274 6040 -4188 6074
rect -4274 6006 -4248 6040
rect -4214 6006 -4188 6040
rect -4274 5972 -4188 6006
rect -4274 5938 -4248 5972
rect -4214 5938 -4188 5972
rect -4274 5884 -4188 5938
rect -3938 6856 -3852 6884
rect -3938 6822 -3912 6856
rect -3878 6822 -3852 6856
rect -3938 6788 -3852 6822
rect -3938 6754 -3912 6788
rect -3878 6754 -3852 6788
rect -3938 6720 -3852 6754
rect -3938 6686 -3912 6720
rect -3878 6686 -3852 6720
rect -3938 6652 -3852 6686
rect -3938 6618 -3912 6652
rect -3878 6618 -3852 6652
rect -3938 6584 -3852 6618
rect -3938 6550 -3912 6584
rect -3878 6550 -3852 6584
rect -3938 6516 -3852 6550
rect -3938 6482 -3912 6516
rect -3878 6482 -3852 6516
rect -3938 6448 -3852 6482
rect -3938 6414 -3912 6448
rect -3878 6414 -3852 6448
rect -3938 6380 -3852 6414
rect -3938 6346 -3912 6380
rect -3878 6346 -3852 6380
rect -3938 6312 -3852 6346
rect -3938 6278 -3912 6312
rect -3878 6278 -3852 6312
rect -3938 6244 -3852 6278
rect -3938 6210 -3912 6244
rect -3878 6210 -3852 6244
rect -3938 6176 -3852 6210
rect -3938 6142 -3912 6176
rect -3878 6142 -3852 6176
rect -3938 6108 -3852 6142
rect -3938 6074 -3912 6108
rect -3878 6074 -3852 6108
rect -3938 6040 -3852 6074
rect -3938 6006 -3912 6040
rect -3878 6006 -3852 6040
rect -3938 5972 -3852 6006
rect -3938 5938 -3912 5972
rect -3878 5938 -3852 5972
rect -3938 5884 -3852 5938
rect -3602 6856 -3516 6884
rect -3602 6822 -3576 6856
rect -3542 6822 -3516 6856
rect -3602 6788 -3516 6822
rect -3602 6754 -3576 6788
rect -3542 6754 -3516 6788
rect -3602 6720 -3516 6754
rect -3602 6686 -3576 6720
rect -3542 6686 -3516 6720
rect -3602 6652 -3516 6686
rect -3602 6618 -3576 6652
rect -3542 6618 -3516 6652
rect -3602 6584 -3516 6618
rect -3602 6550 -3576 6584
rect -3542 6550 -3516 6584
rect -3602 6516 -3516 6550
rect -3602 6482 -3576 6516
rect -3542 6482 -3516 6516
rect -3602 6448 -3516 6482
rect -3602 6414 -3576 6448
rect -3542 6414 -3516 6448
rect -3602 6380 -3516 6414
rect -3602 6346 -3576 6380
rect -3542 6346 -3516 6380
rect -3602 6312 -3516 6346
rect -3602 6278 -3576 6312
rect -3542 6278 -3516 6312
rect -3602 6244 -3516 6278
rect -3602 6210 -3576 6244
rect -3542 6210 -3516 6244
rect -3602 6176 -3516 6210
rect -3602 6142 -3576 6176
rect -3542 6142 -3516 6176
rect -3602 6108 -3516 6142
rect -3602 6074 -3576 6108
rect -3542 6074 -3516 6108
rect -3602 6040 -3516 6074
rect -3602 6006 -3576 6040
rect -3542 6006 -3516 6040
rect -3602 5972 -3516 6006
rect -3602 5938 -3576 5972
rect -3542 5938 -3516 5972
rect -3602 5884 -3516 5938
rect -3266 6856 -3180 6884
rect -3266 6822 -3240 6856
rect -3206 6822 -3180 6856
rect -3266 6788 -3180 6822
rect -3266 6754 -3240 6788
rect -3206 6754 -3180 6788
rect -3266 6720 -3180 6754
rect -3266 6686 -3240 6720
rect -3206 6686 -3180 6720
rect -3266 6652 -3180 6686
rect -3266 6618 -3240 6652
rect -3206 6618 -3180 6652
rect -3266 6584 -3180 6618
rect -3266 6550 -3240 6584
rect -3206 6550 -3180 6584
rect -3266 6516 -3180 6550
rect -3266 6482 -3240 6516
rect -3206 6482 -3180 6516
rect -3266 6448 -3180 6482
rect -3266 6414 -3240 6448
rect -3206 6414 -3180 6448
rect -3266 6380 -3180 6414
rect -3266 6346 -3240 6380
rect -3206 6346 -3180 6380
rect -3266 6312 -3180 6346
rect -3266 6278 -3240 6312
rect -3206 6278 -3180 6312
rect -3266 6244 -3180 6278
rect -3266 6210 -3240 6244
rect -3206 6210 -3180 6244
rect -3266 6176 -3180 6210
rect -3266 6142 -3240 6176
rect -3206 6142 -3180 6176
rect -3266 6108 -3180 6142
rect -3266 6074 -3240 6108
rect -3206 6074 -3180 6108
rect -3266 6040 -3180 6074
rect -3266 6006 -3240 6040
rect -3206 6006 -3180 6040
rect -3266 5972 -3180 6006
rect -3266 5938 -3240 5972
rect -3206 5938 -3180 5972
rect -3266 5884 -3180 5938
rect -2930 6856 -2844 6884
rect -2930 6822 -2904 6856
rect -2870 6822 -2844 6856
rect -2930 6788 -2844 6822
rect -2930 6754 -2904 6788
rect -2870 6754 -2844 6788
rect -2930 6720 -2844 6754
rect -2930 6686 -2904 6720
rect -2870 6686 -2844 6720
rect -2930 6652 -2844 6686
rect -2930 6618 -2904 6652
rect -2870 6618 -2844 6652
rect -2930 6584 -2844 6618
rect -2930 6550 -2904 6584
rect -2870 6550 -2844 6584
rect -2930 6516 -2844 6550
rect -2930 6482 -2904 6516
rect -2870 6482 -2844 6516
rect -2930 6448 -2844 6482
rect -2930 6414 -2904 6448
rect -2870 6414 -2844 6448
rect -2930 6380 -2844 6414
rect -2930 6346 -2904 6380
rect -2870 6346 -2844 6380
rect -2930 6312 -2844 6346
rect -2930 6278 -2904 6312
rect -2870 6278 -2844 6312
rect -2930 6244 -2844 6278
rect -2930 6210 -2904 6244
rect -2870 6210 -2844 6244
rect -2930 6176 -2844 6210
rect -2930 6142 -2904 6176
rect -2870 6142 -2844 6176
rect -2930 6108 -2844 6142
rect -2930 6074 -2904 6108
rect -2870 6074 -2844 6108
rect -2930 6040 -2844 6074
rect -2930 6006 -2904 6040
rect -2870 6006 -2844 6040
rect -2930 5972 -2844 6006
rect -2930 5938 -2904 5972
rect -2870 5938 -2844 5972
rect -2930 5884 -2844 5938
rect -2594 6856 -2530 6884
rect -2594 6822 -2568 6856
rect -2534 6822 -2530 6856
rect -2594 6788 -2530 6822
rect -2594 6754 -2568 6788
rect -2534 6754 -2530 6788
rect -2594 6720 -2530 6754
rect -2594 6686 -2568 6720
rect -2534 6686 -2530 6720
rect -2594 6652 -2530 6686
rect -2594 6618 -2568 6652
rect -2534 6618 -2530 6652
rect -2594 6584 -2530 6618
rect -2594 6550 -2568 6584
rect -2534 6550 -2530 6584
rect -2594 6516 -2530 6550
rect -2594 6482 -2568 6516
rect -2534 6482 -2530 6516
rect -2594 6448 -2530 6482
rect -2594 6414 -2568 6448
rect -2534 6414 -2530 6448
rect -2594 6380 -2530 6414
rect -2594 6346 -2568 6380
rect -2534 6346 -2530 6380
rect -2594 6312 -2530 6346
rect -2594 6278 -2568 6312
rect -2534 6278 -2530 6312
rect -2594 6244 -2530 6278
rect -2594 6210 -2568 6244
rect -2534 6210 -2530 6244
rect -2594 6176 -2530 6210
rect -2594 6142 -2568 6176
rect -2534 6142 -2530 6176
rect -2594 6108 -2530 6142
rect -2594 6074 -2568 6108
rect -2534 6074 -2530 6108
rect -2594 6040 -2530 6074
rect -2594 6006 -2568 6040
rect -2534 6006 -2530 6040
rect -2594 5972 -2530 6006
rect -2594 5938 -2568 5972
rect -2534 5938 -2530 5972
rect -2594 5884 -2530 5938
rect 810 6880 874 6934
rect 810 6846 814 6880
rect 848 6846 874 6880
rect 810 6812 874 6846
rect 810 6778 814 6812
rect 848 6778 874 6812
rect 810 6744 874 6778
rect 810 6710 814 6744
rect 848 6710 874 6744
rect 810 6676 874 6710
rect 810 6642 814 6676
rect 848 6642 874 6676
rect 810 6608 874 6642
rect 810 6574 814 6608
rect 848 6574 874 6608
rect 810 6540 874 6574
rect 810 6506 814 6540
rect 848 6506 874 6540
rect 810 6472 874 6506
rect 810 6438 814 6472
rect 848 6438 874 6472
rect 810 6404 874 6438
rect 810 6370 814 6404
rect 848 6370 874 6404
rect 810 6336 874 6370
rect 810 6302 814 6336
rect 848 6302 874 6336
rect 810 6268 874 6302
rect 810 6234 814 6268
rect 848 6234 874 6268
rect 810 6200 874 6234
rect 810 6166 814 6200
rect 848 6166 874 6200
rect 810 6132 874 6166
rect 810 6098 814 6132
rect 848 6098 874 6132
rect 810 6064 874 6098
rect 810 6030 814 6064
rect 848 6030 874 6064
rect 810 5996 874 6030
rect 810 5962 814 5996
rect 848 5962 874 5996
rect 810 5934 874 5962
rect 1124 6906 1210 6934
rect 1124 6872 1150 6906
rect 1184 6872 1210 6906
rect 1124 6838 1210 6872
rect 1124 6804 1150 6838
rect 1184 6804 1210 6838
rect 1124 6770 1210 6804
rect 1124 6736 1150 6770
rect 1184 6736 1210 6770
rect 1124 6702 1210 6736
rect 1124 6668 1150 6702
rect 1184 6668 1210 6702
rect 1124 6634 1210 6668
rect 1124 6600 1150 6634
rect 1184 6600 1210 6634
rect 1124 6566 1210 6600
rect 1124 6532 1150 6566
rect 1184 6532 1210 6566
rect 1124 6498 1210 6532
rect 1124 6464 1150 6498
rect 1184 6464 1210 6498
rect 1124 6430 1210 6464
rect 1124 6396 1150 6430
rect 1184 6396 1210 6430
rect 1124 6362 1210 6396
rect 1124 6328 1150 6362
rect 1184 6328 1210 6362
rect 1124 6294 1210 6328
rect 1124 6260 1150 6294
rect 1184 6260 1210 6294
rect 1124 6226 1210 6260
rect 1124 6192 1150 6226
rect 1184 6192 1210 6226
rect 1124 6158 1210 6192
rect 1124 6124 1150 6158
rect 1184 6124 1210 6158
rect 1124 6090 1210 6124
rect 1124 6056 1150 6090
rect 1184 6056 1210 6090
rect 1124 6022 1210 6056
rect 1124 5988 1150 6022
rect 1184 5988 1210 6022
rect 1124 5934 1210 5988
rect 1460 6906 1546 6934
rect 1460 6872 1486 6906
rect 1520 6872 1546 6906
rect 1460 6838 1546 6872
rect 1460 6804 1486 6838
rect 1520 6804 1546 6838
rect 1460 6770 1546 6804
rect 1460 6736 1486 6770
rect 1520 6736 1546 6770
rect 1460 6702 1546 6736
rect 1460 6668 1486 6702
rect 1520 6668 1546 6702
rect 1460 6634 1546 6668
rect 1460 6600 1486 6634
rect 1520 6600 1546 6634
rect 1460 6566 1546 6600
rect 1460 6532 1486 6566
rect 1520 6532 1546 6566
rect 1460 6498 1546 6532
rect 1460 6464 1486 6498
rect 1520 6464 1546 6498
rect 1460 6430 1546 6464
rect 1460 6396 1486 6430
rect 1520 6396 1546 6430
rect 1460 6362 1546 6396
rect 1460 6328 1486 6362
rect 1520 6328 1546 6362
rect 1460 6294 1546 6328
rect 1460 6260 1486 6294
rect 1520 6260 1546 6294
rect 1460 6226 1546 6260
rect 1460 6192 1486 6226
rect 1520 6192 1546 6226
rect 1460 6158 1546 6192
rect 1460 6124 1486 6158
rect 1520 6124 1546 6158
rect 1460 6090 1546 6124
rect 1460 6056 1486 6090
rect 1520 6056 1546 6090
rect 1460 6022 1546 6056
rect 1460 5988 1486 6022
rect 1520 5988 1546 6022
rect 1460 5934 1546 5988
rect 1796 6906 1882 6934
rect 1796 6872 1822 6906
rect 1856 6872 1882 6906
rect 1796 6838 1882 6872
rect 1796 6804 1822 6838
rect 1856 6804 1882 6838
rect 1796 6770 1882 6804
rect 1796 6736 1822 6770
rect 1856 6736 1882 6770
rect 1796 6702 1882 6736
rect 1796 6668 1822 6702
rect 1856 6668 1882 6702
rect 1796 6634 1882 6668
rect 1796 6600 1822 6634
rect 1856 6600 1882 6634
rect 1796 6566 1882 6600
rect 1796 6532 1822 6566
rect 1856 6532 1882 6566
rect 1796 6498 1882 6532
rect 1796 6464 1822 6498
rect 1856 6464 1882 6498
rect 1796 6430 1882 6464
rect 1796 6396 1822 6430
rect 1856 6396 1882 6430
rect 1796 6362 1882 6396
rect 1796 6328 1822 6362
rect 1856 6328 1882 6362
rect 1796 6294 1882 6328
rect 1796 6260 1822 6294
rect 1856 6260 1882 6294
rect 1796 6226 1882 6260
rect 1796 6192 1822 6226
rect 1856 6192 1882 6226
rect 1796 6158 1882 6192
rect 1796 6124 1822 6158
rect 1856 6124 1882 6158
rect 1796 6090 1882 6124
rect 1796 6056 1822 6090
rect 1856 6056 1882 6090
rect 1796 6022 1882 6056
rect 1796 5988 1822 6022
rect 1856 5988 1882 6022
rect 1796 5934 1882 5988
rect 2132 6906 2218 6934
rect 2132 6872 2158 6906
rect 2192 6872 2218 6906
rect 2132 6838 2218 6872
rect 2132 6804 2158 6838
rect 2192 6804 2218 6838
rect 2132 6770 2218 6804
rect 2132 6736 2158 6770
rect 2192 6736 2218 6770
rect 2132 6702 2218 6736
rect 2132 6668 2158 6702
rect 2192 6668 2218 6702
rect 2132 6634 2218 6668
rect 2132 6600 2158 6634
rect 2192 6600 2218 6634
rect 2132 6566 2218 6600
rect 2132 6532 2158 6566
rect 2192 6532 2218 6566
rect 2132 6498 2218 6532
rect 2132 6464 2158 6498
rect 2192 6464 2218 6498
rect 2132 6430 2218 6464
rect 2132 6396 2158 6430
rect 2192 6396 2218 6430
rect 2132 6362 2218 6396
rect 2132 6328 2158 6362
rect 2192 6328 2218 6362
rect 2132 6294 2218 6328
rect 2132 6260 2158 6294
rect 2192 6260 2218 6294
rect 2132 6226 2218 6260
rect 2132 6192 2158 6226
rect 2192 6192 2218 6226
rect 2132 6158 2218 6192
rect 2132 6124 2158 6158
rect 2192 6124 2218 6158
rect 2132 6090 2218 6124
rect 2132 6056 2158 6090
rect 2192 6056 2218 6090
rect 2132 6022 2218 6056
rect 2132 5988 2158 6022
rect 2192 5988 2218 6022
rect 2132 5934 2218 5988
rect 2468 6906 2554 6934
rect 2468 6872 2494 6906
rect 2528 6872 2554 6906
rect 2468 6838 2554 6872
rect 2468 6804 2494 6838
rect 2528 6804 2554 6838
rect 2468 6770 2554 6804
rect 2468 6736 2494 6770
rect 2528 6736 2554 6770
rect 2468 6702 2554 6736
rect 2468 6668 2494 6702
rect 2528 6668 2554 6702
rect 2468 6634 2554 6668
rect 2468 6600 2494 6634
rect 2528 6600 2554 6634
rect 2468 6566 2554 6600
rect 2468 6532 2494 6566
rect 2528 6532 2554 6566
rect 2468 6498 2554 6532
rect 2468 6464 2494 6498
rect 2528 6464 2554 6498
rect 2468 6430 2554 6464
rect 2468 6396 2494 6430
rect 2528 6396 2554 6430
rect 2468 6362 2554 6396
rect 2468 6328 2494 6362
rect 2528 6328 2554 6362
rect 2468 6294 2554 6328
rect 2468 6260 2494 6294
rect 2528 6260 2554 6294
rect 2468 6226 2554 6260
rect 2468 6192 2494 6226
rect 2528 6192 2554 6226
rect 2468 6158 2554 6192
rect 2468 6124 2494 6158
rect 2528 6124 2554 6158
rect 2468 6090 2554 6124
rect 2468 6056 2494 6090
rect 2528 6056 2554 6090
rect 2468 6022 2554 6056
rect 2468 5988 2494 6022
rect 2528 5988 2554 6022
rect 2468 5934 2554 5988
rect 2804 6906 2868 6934
rect 2804 6872 2830 6906
rect 2864 6872 2868 6906
rect 2804 6838 2868 6872
rect 2804 6804 2830 6838
rect 2864 6804 2868 6838
rect 2804 6770 2868 6804
rect 2804 6736 2830 6770
rect 2864 6736 2868 6770
rect 2804 6702 2868 6736
rect 2804 6668 2830 6702
rect 2864 6668 2868 6702
rect 2804 6634 2868 6668
rect 2804 6600 2830 6634
rect 2864 6600 2868 6634
rect 2804 6566 2868 6600
rect 2804 6532 2830 6566
rect 2864 6532 2868 6566
rect 2804 6498 2868 6532
rect 2804 6464 2830 6498
rect 2864 6464 2868 6498
rect 2804 6430 2868 6464
rect 2804 6396 2830 6430
rect 2864 6396 2868 6430
rect 2804 6362 2868 6396
rect 2804 6328 2830 6362
rect 2864 6328 2868 6362
rect 2804 6294 2868 6328
rect 2804 6260 2830 6294
rect 2864 6260 2868 6294
rect 2804 6226 2868 6260
rect 2804 6192 2830 6226
rect 2864 6192 2868 6226
rect 2804 6158 2868 6192
rect 2804 6124 2830 6158
rect 2864 6124 2868 6158
rect 2804 6090 2868 6124
rect 2804 6056 2830 6090
rect 2864 6056 2868 6090
rect 2804 6022 2868 6056
rect 2804 5988 2830 6022
rect 2864 5988 2868 6022
rect 2804 5934 2868 5988
rect 7180 6880 7244 6934
rect 7180 6846 7184 6880
rect 7218 6846 7244 6880
rect 7180 6812 7244 6846
rect 7180 6778 7184 6812
rect 7218 6778 7244 6812
rect 7180 6744 7244 6778
rect 7180 6710 7184 6744
rect 7218 6710 7244 6744
rect 7180 6676 7244 6710
rect 7180 6642 7184 6676
rect 7218 6642 7244 6676
rect 7180 6608 7244 6642
rect 7180 6574 7184 6608
rect 7218 6574 7244 6608
rect 7180 6540 7244 6574
rect 7180 6506 7184 6540
rect 7218 6506 7244 6540
rect 7180 6472 7244 6506
rect 7180 6438 7184 6472
rect 7218 6438 7244 6472
rect 7180 6404 7244 6438
rect 7180 6370 7184 6404
rect 7218 6370 7244 6404
rect 7180 6336 7244 6370
rect 7180 6302 7184 6336
rect 7218 6302 7244 6336
rect 7180 6268 7244 6302
rect 7180 6234 7184 6268
rect 7218 6234 7244 6268
rect 7180 6200 7244 6234
rect 7180 6166 7184 6200
rect 7218 6166 7244 6200
rect 7180 6132 7244 6166
rect 7180 6098 7184 6132
rect 7218 6098 7244 6132
rect 7180 6064 7244 6098
rect 7180 6030 7184 6064
rect 7218 6030 7244 6064
rect 7180 5996 7244 6030
rect 7180 5962 7184 5996
rect 7218 5962 7244 5996
rect 7180 5934 7244 5962
rect 7494 6906 7580 6934
rect 7494 6872 7520 6906
rect 7554 6872 7580 6906
rect 7494 6838 7580 6872
rect 7494 6804 7520 6838
rect 7554 6804 7580 6838
rect 7494 6770 7580 6804
rect 7494 6736 7520 6770
rect 7554 6736 7580 6770
rect 7494 6702 7580 6736
rect 7494 6668 7520 6702
rect 7554 6668 7580 6702
rect 7494 6634 7580 6668
rect 7494 6600 7520 6634
rect 7554 6600 7580 6634
rect 7494 6566 7580 6600
rect 7494 6532 7520 6566
rect 7554 6532 7580 6566
rect 7494 6498 7580 6532
rect 7494 6464 7520 6498
rect 7554 6464 7580 6498
rect 7494 6430 7580 6464
rect 7494 6396 7520 6430
rect 7554 6396 7580 6430
rect 7494 6362 7580 6396
rect 7494 6328 7520 6362
rect 7554 6328 7580 6362
rect 7494 6294 7580 6328
rect 7494 6260 7520 6294
rect 7554 6260 7580 6294
rect 7494 6226 7580 6260
rect 7494 6192 7520 6226
rect 7554 6192 7580 6226
rect 7494 6158 7580 6192
rect 7494 6124 7520 6158
rect 7554 6124 7580 6158
rect 7494 6090 7580 6124
rect 7494 6056 7520 6090
rect 7554 6056 7580 6090
rect 7494 6022 7580 6056
rect 7494 5988 7520 6022
rect 7554 5988 7580 6022
rect 7494 5934 7580 5988
rect 7830 6906 7916 6934
rect 7830 6872 7856 6906
rect 7890 6872 7916 6906
rect 7830 6838 7916 6872
rect 7830 6804 7856 6838
rect 7890 6804 7916 6838
rect 7830 6770 7916 6804
rect 7830 6736 7856 6770
rect 7890 6736 7916 6770
rect 7830 6702 7916 6736
rect 7830 6668 7856 6702
rect 7890 6668 7916 6702
rect 7830 6634 7916 6668
rect 7830 6600 7856 6634
rect 7890 6600 7916 6634
rect 7830 6566 7916 6600
rect 7830 6532 7856 6566
rect 7890 6532 7916 6566
rect 7830 6498 7916 6532
rect 7830 6464 7856 6498
rect 7890 6464 7916 6498
rect 7830 6430 7916 6464
rect 7830 6396 7856 6430
rect 7890 6396 7916 6430
rect 7830 6362 7916 6396
rect 7830 6328 7856 6362
rect 7890 6328 7916 6362
rect 7830 6294 7916 6328
rect 7830 6260 7856 6294
rect 7890 6260 7916 6294
rect 7830 6226 7916 6260
rect 7830 6192 7856 6226
rect 7890 6192 7916 6226
rect 7830 6158 7916 6192
rect 7830 6124 7856 6158
rect 7890 6124 7916 6158
rect 7830 6090 7916 6124
rect 7830 6056 7856 6090
rect 7890 6056 7916 6090
rect 7830 6022 7916 6056
rect 7830 5988 7856 6022
rect 7890 5988 7916 6022
rect 7830 5934 7916 5988
rect 8166 6906 8252 6934
rect 8166 6872 8192 6906
rect 8226 6872 8252 6906
rect 8166 6838 8252 6872
rect 8166 6804 8192 6838
rect 8226 6804 8252 6838
rect 8166 6770 8252 6804
rect 8166 6736 8192 6770
rect 8226 6736 8252 6770
rect 8166 6702 8252 6736
rect 8166 6668 8192 6702
rect 8226 6668 8252 6702
rect 8166 6634 8252 6668
rect 8166 6600 8192 6634
rect 8226 6600 8252 6634
rect 8166 6566 8252 6600
rect 8166 6532 8192 6566
rect 8226 6532 8252 6566
rect 8166 6498 8252 6532
rect 8166 6464 8192 6498
rect 8226 6464 8252 6498
rect 8166 6430 8252 6464
rect 8166 6396 8192 6430
rect 8226 6396 8252 6430
rect 8166 6362 8252 6396
rect 8166 6328 8192 6362
rect 8226 6328 8252 6362
rect 8166 6294 8252 6328
rect 8166 6260 8192 6294
rect 8226 6260 8252 6294
rect 8166 6226 8252 6260
rect 8166 6192 8192 6226
rect 8226 6192 8252 6226
rect 8166 6158 8252 6192
rect 8166 6124 8192 6158
rect 8226 6124 8252 6158
rect 8166 6090 8252 6124
rect 8166 6056 8192 6090
rect 8226 6056 8252 6090
rect 8166 6022 8252 6056
rect 8166 5988 8192 6022
rect 8226 5988 8252 6022
rect 8166 5934 8252 5988
rect 8502 6906 8588 6934
rect 8502 6872 8528 6906
rect 8562 6872 8588 6906
rect 8502 6838 8588 6872
rect 8502 6804 8528 6838
rect 8562 6804 8588 6838
rect 8502 6770 8588 6804
rect 8502 6736 8528 6770
rect 8562 6736 8588 6770
rect 8502 6702 8588 6736
rect 8502 6668 8528 6702
rect 8562 6668 8588 6702
rect 8502 6634 8588 6668
rect 8502 6600 8528 6634
rect 8562 6600 8588 6634
rect 8502 6566 8588 6600
rect 8502 6532 8528 6566
rect 8562 6532 8588 6566
rect 8502 6498 8588 6532
rect 8502 6464 8528 6498
rect 8562 6464 8588 6498
rect 8502 6430 8588 6464
rect 8502 6396 8528 6430
rect 8562 6396 8588 6430
rect 8502 6362 8588 6396
rect 8502 6328 8528 6362
rect 8562 6328 8588 6362
rect 8502 6294 8588 6328
rect 8502 6260 8528 6294
rect 8562 6260 8588 6294
rect 8502 6226 8588 6260
rect 8502 6192 8528 6226
rect 8562 6192 8588 6226
rect 8502 6158 8588 6192
rect 8502 6124 8528 6158
rect 8562 6124 8588 6158
rect 8502 6090 8588 6124
rect 8502 6056 8528 6090
rect 8562 6056 8588 6090
rect 8502 6022 8588 6056
rect 8502 5988 8528 6022
rect 8562 5988 8588 6022
rect 8502 5934 8588 5988
rect 8838 6906 8924 6934
rect 8838 6872 8864 6906
rect 8898 6872 8924 6906
rect 8838 6838 8924 6872
rect 8838 6804 8864 6838
rect 8898 6804 8924 6838
rect 8838 6770 8924 6804
rect 8838 6736 8864 6770
rect 8898 6736 8924 6770
rect 8838 6702 8924 6736
rect 8838 6668 8864 6702
rect 8898 6668 8924 6702
rect 8838 6634 8924 6668
rect 8838 6600 8864 6634
rect 8898 6600 8924 6634
rect 8838 6566 8924 6600
rect 8838 6532 8864 6566
rect 8898 6532 8924 6566
rect 8838 6498 8924 6532
rect 8838 6464 8864 6498
rect 8898 6464 8924 6498
rect 8838 6430 8924 6464
rect 8838 6396 8864 6430
rect 8898 6396 8924 6430
rect 8838 6362 8924 6396
rect 8838 6328 8864 6362
rect 8898 6328 8924 6362
rect 8838 6294 8924 6328
rect 8838 6260 8864 6294
rect 8898 6260 8924 6294
rect 8838 6226 8924 6260
rect 8838 6192 8864 6226
rect 8898 6192 8924 6226
rect 8838 6158 8924 6192
rect 8838 6124 8864 6158
rect 8898 6124 8924 6158
rect 8838 6090 8924 6124
rect 8838 6056 8864 6090
rect 8898 6056 8924 6090
rect 8838 6022 8924 6056
rect 8838 5988 8864 6022
rect 8898 5988 8924 6022
rect 8838 5934 8924 5988
rect 9174 6906 9238 6934
rect 9174 6872 9200 6906
rect 9234 6872 9238 6906
rect 9174 6838 9238 6872
rect 9174 6804 9200 6838
rect 9234 6804 9238 6838
rect 9174 6770 9238 6804
rect 9174 6736 9200 6770
rect 9234 6736 9238 6770
rect 9174 6702 9238 6736
rect 9174 6668 9200 6702
rect 9234 6668 9238 6702
rect 9174 6634 9238 6668
rect 9174 6600 9200 6634
rect 9234 6600 9238 6634
rect 9174 6566 9238 6600
rect 9174 6532 9200 6566
rect 9234 6532 9238 6566
rect 9174 6498 9238 6532
rect 9174 6464 9200 6498
rect 9234 6464 9238 6498
rect 9174 6430 9238 6464
rect 9174 6396 9200 6430
rect 9234 6396 9238 6430
rect 9174 6362 9238 6396
rect 9174 6328 9200 6362
rect 9234 6328 9238 6362
rect 9174 6294 9238 6328
rect 9174 6260 9200 6294
rect 9234 6260 9238 6294
rect 9174 6226 9238 6260
rect 9174 6192 9200 6226
rect 9234 6192 9238 6226
rect 9174 6158 9238 6192
rect 9174 6124 9200 6158
rect 9234 6124 9238 6158
rect 9174 6090 9238 6124
rect 9174 6056 9200 6090
rect 9234 6056 9238 6090
rect 9174 6022 9238 6056
rect 9174 5988 9200 6022
rect 9234 5988 9238 6022
rect 9174 5934 9238 5988
rect 13550 6880 13614 6934
rect 13550 6846 13554 6880
rect 13588 6846 13614 6880
rect 13550 6812 13614 6846
rect 13550 6778 13554 6812
rect 13588 6778 13614 6812
rect 13550 6744 13614 6778
rect 13550 6710 13554 6744
rect 13588 6710 13614 6744
rect 13550 6676 13614 6710
rect 13550 6642 13554 6676
rect 13588 6642 13614 6676
rect 13550 6608 13614 6642
rect 13550 6574 13554 6608
rect 13588 6574 13614 6608
rect 13550 6540 13614 6574
rect 13550 6506 13554 6540
rect 13588 6506 13614 6540
rect 13550 6472 13614 6506
rect 13550 6438 13554 6472
rect 13588 6438 13614 6472
rect 13550 6404 13614 6438
rect 13550 6370 13554 6404
rect 13588 6370 13614 6404
rect 13550 6336 13614 6370
rect 13550 6302 13554 6336
rect 13588 6302 13614 6336
rect 13550 6268 13614 6302
rect 13550 6234 13554 6268
rect 13588 6234 13614 6268
rect 13550 6200 13614 6234
rect 13550 6166 13554 6200
rect 13588 6166 13614 6200
rect 13550 6132 13614 6166
rect 13550 6098 13554 6132
rect 13588 6098 13614 6132
rect 13550 6064 13614 6098
rect 13550 6030 13554 6064
rect 13588 6030 13614 6064
rect 13550 5996 13614 6030
rect 13550 5962 13554 5996
rect 13588 5962 13614 5996
rect 13550 5934 13614 5962
rect 13864 6906 13950 6934
rect 13864 6872 13890 6906
rect 13924 6872 13950 6906
rect 13864 6838 13950 6872
rect 13864 6804 13890 6838
rect 13924 6804 13950 6838
rect 13864 6770 13950 6804
rect 13864 6736 13890 6770
rect 13924 6736 13950 6770
rect 13864 6702 13950 6736
rect 13864 6668 13890 6702
rect 13924 6668 13950 6702
rect 13864 6634 13950 6668
rect 13864 6600 13890 6634
rect 13924 6600 13950 6634
rect 13864 6566 13950 6600
rect 13864 6532 13890 6566
rect 13924 6532 13950 6566
rect 13864 6498 13950 6532
rect 13864 6464 13890 6498
rect 13924 6464 13950 6498
rect 13864 6430 13950 6464
rect 13864 6396 13890 6430
rect 13924 6396 13950 6430
rect 13864 6362 13950 6396
rect 13864 6328 13890 6362
rect 13924 6328 13950 6362
rect 13864 6294 13950 6328
rect 13864 6260 13890 6294
rect 13924 6260 13950 6294
rect 13864 6226 13950 6260
rect 13864 6192 13890 6226
rect 13924 6192 13950 6226
rect 13864 6158 13950 6192
rect 13864 6124 13890 6158
rect 13924 6124 13950 6158
rect 13864 6090 13950 6124
rect 13864 6056 13890 6090
rect 13924 6056 13950 6090
rect 13864 6022 13950 6056
rect 13864 5988 13890 6022
rect 13924 5988 13950 6022
rect 13864 5934 13950 5988
rect 14200 6906 14286 6934
rect 14200 6872 14226 6906
rect 14260 6872 14286 6906
rect 14200 6838 14286 6872
rect 14200 6804 14226 6838
rect 14260 6804 14286 6838
rect 14200 6770 14286 6804
rect 14200 6736 14226 6770
rect 14260 6736 14286 6770
rect 14200 6702 14286 6736
rect 14200 6668 14226 6702
rect 14260 6668 14286 6702
rect 14200 6634 14286 6668
rect 14200 6600 14226 6634
rect 14260 6600 14286 6634
rect 14200 6566 14286 6600
rect 14200 6532 14226 6566
rect 14260 6532 14286 6566
rect 14200 6498 14286 6532
rect 14200 6464 14226 6498
rect 14260 6464 14286 6498
rect 14200 6430 14286 6464
rect 14200 6396 14226 6430
rect 14260 6396 14286 6430
rect 14200 6362 14286 6396
rect 14200 6328 14226 6362
rect 14260 6328 14286 6362
rect 14200 6294 14286 6328
rect 14200 6260 14226 6294
rect 14260 6260 14286 6294
rect 14200 6226 14286 6260
rect 14200 6192 14226 6226
rect 14260 6192 14286 6226
rect 14200 6158 14286 6192
rect 14200 6124 14226 6158
rect 14260 6124 14286 6158
rect 14200 6090 14286 6124
rect 14200 6056 14226 6090
rect 14260 6056 14286 6090
rect 14200 6022 14286 6056
rect 14200 5988 14226 6022
rect 14260 5988 14286 6022
rect 14200 5934 14286 5988
rect 14536 6906 14622 6934
rect 14536 6872 14562 6906
rect 14596 6872 14622 6906
rect 14536 6838 14622 6872
rect 14536 6804 14562 6838
rect 14596 6804 14622 6838
rect 14536 6770 14622 6804
rect 14536 6736 14562 6770
rect 14596 6736 14622 6770
rect 14536 6702 14622 6736
rect 14536 6668 14562 6702
rect 14596 6668 14622 6702
rect 14536 6634 14622 6668
rect 14536 6600 14562 6634
rect 14596 6600 14622 6634
rect 14536 6566 14622 6600
rect 14536 6532 14562 6566
rect 14596 6532 14622 6566
rect 14536 6498 14622 6532
rect 14536 6464 14562 6498
rect 14596 6464 14622 6498
rect 14536 6430 14622 6464
rect 14536 6396 14562 6430
rect 14596 6396 14622 6430
rect 14536 6362 14622 6396
rect 14536 6328 14562 6362
rect 14596 6328 14622 6362
rect 14536 6294 14622 6328
rect 14536 6260 14562 6294
rect 14596 6260 14622 6294
rect 14536 6226 14622 6260
rect 14536 6192 14562 6226
rect 14596 6192 14622 6226
rect 14536 6158 14622 6192
rect 14536 6124 14562 6158
rect 14596 6124 14622 6158
rect 14536 6090 14622 6124
rect 14536 6056 14562 6090
rect 14596 6056 14622 6090
rect 14536 6022 14622 6056
rect 14536 5988 14562 6022
rect 14596 5988 14622 6022
rect 14536 5934 14622 5988
rect 14872 6906 14958 6934
rect 14872 6872 14898 6906
rect 14932 6872 14958 6906
rect 14872 6838 14958 6872
rect 14872 6804 14898 6838
rect 14932 6804 14958 6838
rect 14872 6770 14958 6804
rect 14872 6736 14898 6770
rect 14932 6736 14958 6770
rect 14872 6702 14958 6736
rect 14872 6668 14898 6702
rect 14932 6668 14958 6702
rect 14872 6634 14958 6668
rect 14872 6600 14898 6634
rect 14932 6600 14958 6634
rect 14872 6566 14958 6600
rect 14872 6532 14898 6566
rect 14932 6532 14958 6566
rect 14872 6498 14958 6532
rect 14872 6464 14898 6498
rect 14932 6464 14958 6498
rect 14872 6430 14958 6464
rect 14872 6396 14898 6430
rect 14932 6396 14958 6430
rect 14872 6362 14958 6396
rect 14872 6328 14898 6362
rect 14932 6328 14958 6362
rect 14872 6294 14958 6328
rect 14872 6260 14898 6294
rect 14932 6260 14958 6294
rect 14872 6226 14958 6260
rect 14872 6192 14898 6226
rect 14932 6192 14958 6226
rect 14872 6158 14958 6192
rect 14872 6124 14898 6158
rect 14932 6124 14958 6158
rect 14872 6090 14958 6124
rect 14872 6056 14898 6090
rect 14932 6056 14958 6090
rect 14872 6022 14958 6056
rect 14872 5988 14898 6022
rect 14932 5988 14958 6022
rect 14872 5934 14958 5988
rect 15208 6906 15294 6934
rect 15208 6872 15234 6906
rect 15268 6872 15294 6906
rect 15208 6838 15294 6872
rect 15208 6804 15234 6838
rect 15268 6804 15294 6838
rect 15208 6770 15294 6804
rect 15208 6736 15234 6770
rect 15268 6736 15294 6770
rect 15208 6702 15294 6736
rect 15208 6668 15234 6702
rect 15268 6668 15294 6702
rect 15208 6634 15294 6668
rect 15208 6600 15234 6634
rect 15268 6600 15294 6634
rect 15208 6566 15294 6600
rect 15208 6532 15234 6566
rect 15268 6532 15294 6566
rect 15208 6498 15294 6532
rect 15208 6464 15234 6498
rect 15268 6464 15294 6498
rect 15208 6430 15294 6464
rect 15208 6396 15234 6430
rect 15268 6396 15294 6430
rect 15208 6362 15294 6396
rect 15208 6328 15234 6362
rect 15268 6328 15294 6362
rect 15208 6294 15294 6328
rect 15208 6260 15234 6294
rect 15268 6260 15294 6294
rect 15208 6226 15294 6260
rect 15208 6192 15234 6226
rect 15268 6192 15294 6226
rect 15208 6158 15294 6192
rect 15208 6124 15234 6158
rect 15268 6124 15294 6158
rect 15208 6090 15294 6124
rect 15208 6056 15234 6090
rect 15268 6056 15294 6090
rect 15208 6022 15294 6056
rect 15208 5988 15234 6022
rect 15268 5988 15294 6022
rect 15208 5934 15294 5988
rect 15544 6906 15608 6934
rect 15544 6872 15570 6906
rect 15604 6872 15608 6906
rect 15544 6838 15608 6872
rect 15544 6804 15570 6838
rect 15604 6804 15608 6838
rect 15544 6770 15608 6804
rect 15544 6736 15570 6770
rect 15604 6736 15608 6770
rect 15544 6702 15608 6736
rect 15544 6668 15570 6702
rect 15604 6668 15608 6702
rect 15544 6634 15608 6668
rect 15544 6600 15570 6634
rect 15604 6600 15608 6634
rect 15544 6566 15608 6600
rect 15544 6532 15570 6566
rect 15604 6532 15608 6566
rect 15544 6498 15608 6532
rect 15544 6464 15570 6498
rect 15604 6464 15608 6498
rect 15544 6430 15608 6464
rect 15544 6396 15570 6430
rect 15604 6396 15608 6430
rect 15544 6362 15608 6396
rect 15544 6328 15570 6362
rect 15604 6328 15608 6362
rect 15544 6294 15608 6328
rect 15544 6260 15570 6294
rect 15604 6260 15608 6294
rect 15544 6226 15608 6260
rect 15544 6192 15570 6226
rect 15604 6192 15608 6226
rect 15544 6158 15608 6192
rect 15544 6124 15570 6158
rect 15604 6124 15608 6158
rect 15544 6090 15608 6124
rect 15544 6056 15570 6090
rect 15604 6056 15608 6090
rect 15544 6022 15608 6056
rect 15544 5988 15570 6022
rect 15604 5988 15608 6022
rect 15544 5934 15608 5988
rect 19920 6880 19984 6934
rect 19920 6846 19924 6880
rect 19958 6846 19984 6880
rect 19920 6812 19984 6846
rect 19920 6778 19924 6812
rect 19958 6778 19984 6812
rect 19920 6744 19984 6778
rect 19920 6710 19924 6744
rect 19958 6710 19984 6744
rect 19920 6676 19984 6710
rect 19920 6642 19924 6676
rect 19958 6642 19984 6676
rect 19920 6608 19984 6642
rect 19920 6574 19924 6608
rect 19958 6574 19984 6608
rect 19920 6540 19984 6574
rect 19920 6506 19924 6540
rect 19958 6506 19984 6540
rect 19920 6472 19984 6506
rect 19920 6438 19924 6472
rect 19958 6438 19984 6472
rect 19920 6404 19984 6438
rect 19920 6370 19924 6404
rect 19958 6370 19984 6404
rect 19920 6336 19984 6370
rect 19920 6302 19924 6336
rect 19958 6302 19984 6336
rect 19920 6268 19984 6302
rect 19920 6234 19924 6268
rect 19958 6234 19984 6268
rect 19920 6200 19984 6234
rect 19920 6166 19924 6200
rect 19958 6166 19984 6200
rect 19920 6132 19984 6166
rect 19920 6098 19924 6132
rect 19958 6098 19984 6132
rect 19920 6064 19984 6098
rect 19920 6030 19924 6064
rect 19958 6030 19984 6064
rect 19920 5996 19984 6030
rect 19920 5962 19924 5996
rect 19958 5962 19984 5996
rect 19920 5934 19984 5962
rect 20234 6906 20320 6934
rect 20234 6872 20260 6906
rect 20294 6872 20320 6906
rect 20234 6838 20320 6872
rect 20234 6804 20260 6838
rect 20294 6804 20320 6838
rect 20234 6770 20320 6804
rect 20234 6736 20260 6770
rect 20294 6736 20320 6770
rect 20234 6702 20320 6736
rect 20234 6668 20260 6702
rect 20294 6668 20320 6702
rect 20234 6634 20320 6668
rect 20234 6600 20260 6634
rect 20294 6600 20320 6634
rect 20234 6566 20320 6600
rect 20234 6532 20260 6566
rect 20294 6532 20320 6566
rect 20234 6498 20320 6532
rect 20234 6464 20260 6498
rect 20294 6464 20320 6498
rect 20234 6430 20320 6464
rect 20234 6396 20260 6430
rect 20294 6396 20320 6430
rect 20234 6362 20320 6396
rect 20234 6328 20260 6362
rect 20294 6328 20320 6362
rect 20234 6294 20320 6328
rect 20234 6260 20260 6294
rect 20294 6260 20320 6294
rect 20234 6226 20320 6260
rect 20234 6192 20260 6226
rect 20294 6192 20320 6226
rect 20234 6158 20320 6192
rect 20234 6124 20260 6158
rect 20294 6124 20320 6158
rect 20234 6090 20320 6124
rect 20234 6056 20260 6090
rect 20294 6056 20320 6090
rect 20234 6022 20320 6056
rect 20234 5988 20260 6022
rect 20294 5988 20320 6022
rect 20234 5934 20320 5988
rect 20570 6906 20656 6934
rect 20570 6872 20596 6906
rect 20630 6872 20656 6906
rect 20570 6838 20656 6872
rect 20570 6804 20596 6838
rect 20630 6804 20656 6838
rect 20570 6770 20656 6804
rect 20570 6736 20596 6770
rect 20630 6736 20656 6770
rect 20570 6702 20656 6736
rect 20570 6668 20596 6702
rect 20630 6668 20656 6702
rect 20570 6634 20656 6668
rect 20570 6600 20596 6634
rect 20630 6600 20656 6634
rect 20570 6566 20656 6600
rect 20570 6532 20596 6566
rect 20630 6532 20656 6566
rect 20570 6498 20656 6532
rect 20570 6464 20596 6498
rect 20630 6464 20656 6498
rect 20570 6430 20656 6464
rect 20570 6396 20596 6430
rect 20630 6396 20656 6430
rect 20570 6362 20656 6396
rect 20570 6328 20596 6362
rect 20630 6328 20656 6362
rect 20570 6294 20656 6328
rect 20570 6260 20596 6294
rect 20630 6260 20656 6294
rect 20570 6226 20656 6260
rect 20570 6192 20596 6226
rect 20630 6192 20656 6226
rect 20570 6158 20656 6192
rect 20570 6124 20596 6158
rect 20630 6124 20656 6158
rect 20570 6090 20656 6124
rect 20570 6056 20596 6090
rect 20630 6056 20656 6090
rect 20570 6022 20656 6056
rect 20570 5988 20596 6022
rect 20630 5988 20656 6022
rect 20570 5934 20656 5988
rect 20906 6906 20992 6934
rect 20906 6872 20932 6906
rect 20966 6872 20992 6906
rect 20906 6838 20992 6872
rect 20906 6804 20932 6838
rect 20966 6804 20992 6838
rect 20906 6770 20992 6804
rect 20906 6736 20932 6770
rect 20966 6736 20992 6770
rect 20906 6702 20992 6736
rect 20906 6668 20932 6702
rect 20966 6668 20992 6702
rect 20906 6634 20992 6668
rect 20906 6600 20932 6634
rect 20966 6600 20992 6634
rect 20906 6566 20992 6600
rect 20906 6532 20932 6566
rect 20966 6532 20992 6566
rect 20906 6498 20992 6532
rect 20906 6464 20932 6498
rect 20966 6464 20992 6498
rect 20906 6430 20992 6464
rect 20906 6396 20932 6430
rect 20966 6396 20992 6430
rect 20906 6362 20992 6396
rect 20906 6328 20932 6362
rect 20966 6328 20992 6362
rect 20906 6294 20992 6328
rect 20906 6260 20932 6294
rect 20966 6260 20992 6294
rect 20906 6226 20992 6260
rect 20906 6192 20932 6226
rect 20966 6192 20992 6226
rect 20906 6158 20992 6192
rect 20906 6124 20932 6158
rect 20966 6124 20992 6158
rect 20906 6090 20992 6124
rect 20906 6056 20932 6090
rect 20966 6056 20992 6090
rect 20906 6022 20992 6056
rect 20906 5988 20932 6022
rect 20966 5988 20992 6022
rect 20906 5934 20992 5988
rect 21242 6906 21328 6934
rect 21242 6872 21268 6906
rect 21302 6872 21328 6906
rect 21242 6838 21328 6872
rect 21242 6804 21268 6838
rect 21302 6804 21328 6838
rect 21242 6770 21328 6804
rect 21242 6736 21268 6770
rect 21302 6736 21328 6770
rect 21242 6702 21328 6736
rect 21242 6668 21268 6702
rect 21302 6668 21328 6702
rect 21242 6634 21328 6668
rect 21242 6600 21268 6634
rect 21302 6600 21328 6634
rect 21242 6566 21328 6600
rect 21242 6532 21268 6566
rect 21302 6532 21328 6566
rect 21242 6498 21328 6532
rect 21242 6464 21268 6498
rect 21302 6464 21328 6498
rect 21242 6430 21328 6464
rect 21242 6396 21268 6430
rect 21302 6396 21328 6430
rect 21242 6362 21328 6396
rect 21242 6328 21268 6362
rect 21302 6328 21328 6362
rect 21242 6294 21328 6328
rect 21242 6260 21268 6294
rect 21302 6260 21328 6294
rect 21242 6226 21328 6260
rect 21242 6192 21268 6226
rect 21302 6192 21328 6226
rect 21242 6158 21328 6192
rect 21242 6124 21268 6158
rect 21302 6124 21328 6158
rect 21242 6090 21328 6124
rect 21242 6056 21268 6090
rect 21302 6056 21328 6090
rect 21242 6022 21328 6056
rect 21242 5988 21268 6022
rect 21302 5988 21328 6022
rect 21242 5934 21328 5988
rect 21578 6906 21664 6934
rect 21578 6872 21604 6906
rect 21638 6872 21664 6906
rect 21578 6838 21664 6872
rect 21578 6804 21604 6838
rect 21638 6804 21664 6838
rect 21578 6770 21664 6804
rect 21578 6736 21604 6770
rect 21638 6736 21664 6770
rect 21578 6702 21664 6736
rect 21578 6668 21604 6702
rect 21638 6668 21664 6702
rect 21578 6634 21664 6668
rect 21578 6600 21604 6634
rect 21638 6600 21664 6634
rect 21578 6566 21664 6600
rect 21578 6532 21604 6566
rect 21638 6532 21664 6566
rect 21578 6498 21664 6532
rect 21578 6464 21604 6498
rect 21638 6464 21664 6498
rect 21578 6430 21664 6464
rect 21578 6396 21604 6430
rect 21638 6396 21664 6430
rect 21578 6362 21664 6396
rect 21578 6328 21604 6362
rect 21638 6328 21664 6362
rect 21578 6294 21664 6328
rect 21578 6260 21604 6294
rect 21638 6260 21664 6294
rect 21578 6226 21664 6260
rect 21578 6192 21604 6226
rect 21638 6192 21664 6226
rect 21578 6158 21664 6192
rect 21578 6124 21604 6158
rect 21638 6124 21664 6158
rect 21578 6090 21664 6124
rect 21578 6056 21604 6090
rect 21638 6056 21664 6090
rect 21578 6022 21664 6056
rect 21578 5988 21604 6022
rect 21638 5988 21664 6022
rect 21578 5934 21664 5988
rect 21914 6906 21978 6934
rect 21914 6872 21940 6906
rect 21974 6872 21978 6906
rect 21914 6838 21978 6872
rect 21914 6804 21940 6838
rect 21974 6804 21978 6838
rect 21914 6770 21978 6804
rect 21914 6736 21940 6770
rect 21974 6736 21978 6770
rect 21914 6702 21978 6736
rect 21914 6668 21940 6702
rect 21974 6668 21978 6702
rect 21914 6634 21978 6668
rect 21914 6600 21940 6634
rect 21974 6600 21978 6634
rect 21914 6566 21978 6600
rect 21914 6532 21940 6566
rect 21974 6532 21978 6566
rect 21914 6498 21978 6532
rect 21914 6464 21940 6498
rect 21974 6464 21978 6498
rect 21914 6430 21978 6464
rect 21914 6396 21940 6430
rect 21974 6396 21978 6430
rect 21914 6362 21978 6396
rect 21914 6328 21940 6362
rect 21974 6328 21978 6362
rect 21914 6294 21978 6328
rect 21914 6260 21940 6294
rect 21974 6260 21978 6294
rect 21914 6226 21978 6260
rect 21914 6192 21940 6226
rect 21974 6192 21978 6226
rect 21914 6158 21978 6192
rect 21914 6124 21940 6158
rect 21974 6124 21978 6158
rect 21914 6090 21978 6124
rect 21914 6056 21940 6090
rect 21974 6056 21978 6090
rect 21914 6022 21978 6056
rect 21914 5988 21940 6022
rect 21974 5988 21978 6022
rect 21914 5934 21978 5988
rect 29178 6880 29242 6934
rect 29178 6846 29182 6880
rect 29216 6846 29242 6880
rect 29178 6812 29242 6846
rect 29178 6778 29182 6812
rect 29216 6778 29242 6812
rect 29178 6744 29242 6778
rect 29178 6710 29182 6744
rect 29216 6710 29242 6744
rect 29178 6676 29242 6710
rect 29178 6642 29182 6676
rect 29216 6642 29242 6676
rect 29178 6608 29242 6642
rect 29178 6574 29182 6608
rect 29216 6574 29242 6608
rect 29178 6540 29242 6574
rect 29178 6506 29182 6540
rect 29216 6506 29242 6540
rect 29178 6472 29242 6506
rect 29178 6438 29182 6472
rect 29216 6438 29242 6472
rect 29178 6404 29242 6438
rect 29178 6370 29182 6404
rect 29216 6370 29242 6404
rect 29178 6336 29242 6370
rect 29178 6302 29182 6336
rect 29216 6302 29242 6336
rect 29178 6268 29242 6302
rect 29178 6234 29182 6268
rect 29216 6234 29242 6268
rect 29178 6200 29242 6234
rect 29178 6166 29182 6200
rect 29216 6166 29242 6200
rect 29178 6132 29242 6166
rect 29178 6098 29182 6132
rect 29216 6098 29242 6132
rect 29178 6064 29242 6098
rect 29178 6030 29182 6064
rect 29216 6030 29242 6064
rect 29178 5996 29242 6030
rect 29178 5962 29182 5996
rect 29216 5962 29242 5996
rect 29178 5934 29242 5962
rect 29492 6906 29578 6934
rect 29492 6872 29518 6906
rect 29552 6872 29578 6906
rect 29492 6838 29578 6872
rect 29492 6804 29518 6838
rect 29552 6804 29578 6838
rect 29492 6770 29578 6804
rect 29492 6736 29518 6770
rect 29552 6736 29578 6770
rect 29492 6702 29578 6736
rect 29492 6668 29518 6702
rect 29552 6668 29578 6702
rect 29492 6634 29578 6668
rect 29492 6600 29518 6634
rect 29552 6600 29578 6634
rect 29492 6566 29578 6600
rect 29492 6532 29518 6566
rect 29552 6532 29578 6566
rect 29492 6498 29578 6532
rect 29492 6464 29518 6498
rect 29552 6464 29578 6498
rect 29492 6430 29578 6464
rect 29492 6396 29518 6430
rect 29552 6396 29578 6430
rect 29492 6362 29578 6396
rect 29492 6328 29518 6362
rect 29552 6328 29578 6362
rect 29492 6294 29578 6328
rect 29492 6260 29518 6294
rect 29552 6260 29578 6294
rect 29492 6226 29578 6260
rect 29492 6192 29518 6226
rect 29552 6192 29578 6226
rect 29492 6158 29578 6192
rect 29492 6124 29518 6158
rect 29552 6124 29578 6158
rect 29492 6090 29578 6124
rect 29492 6056 29518 6090
rect 29552 6056 29578 6090
rect 29492 6022 29578 6056
rect 29492 5988 29518 6022
rect 29552 5988 29578 6022
rect 29492 5934 29578 5988
rect 29828 6906 29914 6934
rect 29828 6872 29854 6906
rect 29888 6872 29914 6906
rect 29828 6838 29914 6872
rect 29828 6804 29854 6838
rect 29888 6804 29914 6838
rect 29828 6770 29914 6804
rect 29828 6736 29854 6770
rect 29888 6736 29914 6770
rect 29828 6702 29914 6736
rect 29828 6668 29854 6702
rect 29888 6668 29914 6702
rect 29828 6634 29914 6668
rect 29828 6600 29854 6634
rect 29888 6600 29914 6634
rect 29828 6566 29914 6600
rect 29828 6532 29854 6566
rect 29888 6532 29914 6566
rect 29828 6498 29914 6532
rect 29828 6464 29854 6498
rect 29888 6464 29914 6498
rect 29828 6430 29914 6464
rect 29828 6396 29854 6430
rect 29888 6396 29914 6430
rect 29828 6362 29914 6396
rect 29828 6328 29854 6362
rect 29888 6328 29914 6362
rect 29828 6294 29914 6328
rect 29828 6260 29854 6294
rect 29888 6260 29914 6294
rect 29828 6226 29914 6260
rect 29828 6192 29854 6226
rect 29888 6192 29914 6226
rect 29828 6158 29914 6192
rect 29828 6124 29854 6158
rect 29888 6124 29914 6158
rect 29828 6090 29914 6124
rect 29828 6056 29854 6090
rect 29888 6056 29914 6090
rect 29828 6022 29914 6056
rect 29828 5988 29854 6022
rect 29888 5988 29914 6022
rect 29828 5934 29914 5988
rect 30164 6906 30250 6934
rect 30164 6872 30190 6906
rect 30224 6872 30250 6906
rect 30164 6838 30250 6872
rect 30164 6804 30190 6838
rect 30224 6804 30250 6838
rect 30164 6770 30250 6804
rect 30164 6736 30190 6770
rect 30224 6736 30250 6770
rect 30164 6702 30250 6736
rect 30164 6668 30190 6702
rect 30224 6668 30250 6702
rect 30164 6634 30250 6668
rect 30164 6600 30190 6634
rect 30224 6600 30250 6634
rect 30164 6566 30250 6600
rect 30164 6532 30190 6566
rect 30224 6532 30250 6566
rect 30164 6498 30250 6532
rect 30164 6464 30190 6498
rect 30224 6464 30250 6498
rect 30164 6430 30250 6464
rect 30164 6396 30190 6430
rect 30224 6396 30250 6430
rect 30164 6362 30250 6396
rect 30164 6328 30190 6362
rect 30224 6328 30250 6362
rect 30164 6294 30250 6328
rect 30164 6260 30190 6294
rect 30224 6260 30250 6294
rect 30164 6226 30250 6260
rect 30164 6192 30190 6226
rect 30224 6192 30250 6226
rect 30164 6158 30250 6192
rect 30164 6124 30190 6158
rect 30224 6124 30250 6158
rect 30164 6090 30250 6124
rect 30164 6056 30190 6090
rect 30224 6056 30250 6090
rect 30164 6022 30250 6056
rect 30164 5988 30190 6022
rect 30224 5988 30250 6022
rect 30164 5934 30250 5988
rect 30500 6906 30586 6934
rect 30500 6872 30526 6906
rect 30560 6872 30586 6906
rect 30500 6838 30586 6872
rect 30500 6804 30526 6838
rect 30560 6804 30586 6838
rect 30500 6770 30586 6804
rect 30500 6736 30526 6770
rect 30560 6736 30586 6770
rect 30500 6702 30586 6736
rect 30500 6668 30526 6702
rect 30560 6668 30586 6702
rect 30500 6634 30586 6668
rect 30500 6600 30526 6634
rect 30560 6600 30586 6634
rect 30500 6566 30586 6600
rect 30500 6532 30526 6566
rect 30560 6532 30586 6566
rect 30500 6498 30586 6532
rect 30500 6464 30526 6498
rect 30560 6464 30586 6498
rect 30500 6430 30586 6464
rect 30500 6396 30526 6430
rect 30560 6396 30586 6430
rect 30500 6362 30586 6396
rect 30500 6328 30526 6362
rect 30560 6328 30586 6362
rect 30500 6294 30586 6328
rect 30500 6260 30526 6294
rect 30560 6260 30586 6294
rect 30500 6226 30586 6260
rect 30500 6192 30526 6226
rect 30560 6192 30586 6226
rect 30500 6158 30586 6192
rect 30500 6124 30526 6158
rect 30560 6124 30586 6158
rect 30500 6090 30586 6124
rect 30500 6056 30526 6090
rect 30560 6056 30586 6090
rect 30500 6022 30586 6056
rect 30500 5988 30526 6022
rect 30560 5988 30586 6022
rect 30500 5934 30586 5988
rect 30836 6906 30922 6934
rect 30836 6872 30862 6906
rect 30896 6872 30922 6906
rect 30836 6838 30922 6872
rect 30836 6804 30862 6838
rect 30896 6804 30922 6838
rect 30836 6770 30922 6804
rect 30836 6736 30862 6770
rect 30896 6736 30922 6770
rect 30836 6702 30922 6736
rect 30836 6668 30862 6702
rect 30896 6668 30922 6702
rect 30836 6634 30922 6668
rect 30836 6600 30862 6634
rect 30896 6600 30922 6634
rect 30836 6566 30922 6600
rect 30836 6532 30862 6566
rect 30896 6532 30922 6566
rect 30836 6498 30922 6532
rect 30836 6464 30862 6498
rect 30896 6464 30922 6498
rect 30836 6430 30922 6464
rect 30836 6396 30862 6430
rect 30896 6396 30922 6430
rect 30836 6362 30922 6396
rect 30836 6328 30862 6362
rect 30896 6328 30922 6362
rect 30836 6294 30922 6328
rect 30836 6260 30862 6294
rect 30896 6260 30922 6294
rect 30836 6226 30922 6260
rect 30836 6192 30862 6226
rect 30896 6192 30922 6226
rect 30836 6158 30922 6192
rect 30836 6124 30862 6158
rect 30896 6124 30922 6158
rect 30836 6090 30922 6124
rect 30836 6056 30862 6090
rect 30896 6056 30922 6090
rect 30836 6022 30922 6056
rect 30836 5988 30862 6022
rect 30896 5988 30922 6022
rect 30836 5934 30922 5988
rect 31172 6906 31236 6934
rect 31172 6872 31198 6906
rect 31232 6872 31236 6906
rect 31172 6838 31236 6872
rect 31172 6804 31198 6838
rect 31232 6804 31236 6838
rect 31172 6770 31236 6804
rect 31172 6736 31198 6770
rect 31232 6736 31236 6770
rect 31172 6702 31236 6736
rect 31172 6668 31198 6702
rect 31232 6668 31236 6702
rect 31172 6634 31236 6668
rect 31172 6600 31198 6634
rect 31232 6600 31236 6634
rect 31172 6566 31236 6600
rect 31172 6532 31198 6566
rect 31232 6532 31236 6566
rect 31172 6498 31236 6532
rect 31172 6464 31198 6498
rect 31232 6464 31236 6498
rect 31172 6430 31236 6464
rect 31172 6396 31198 6430
rect 31232 6396 31236 6430
rect 31172 6362 31236 6396
rect 31172 6328 31198 6362
rect 31232 6328 31236 6362
rect 31172 6294 31236 6328
rect 31172 6260 31198 6294
rect 31232 6260 31236 6294
rect 31172 6226 31236 6260
rect 31172 6192 31198 6226
rect 31232 6192 31236 6226
rect 31172 6158 31236 6192
rect 31172 6124 31198 6158
rect 31232 6124 31236 6158
rect 31172 6090 31236 6124
rect 31172 6056 31198 6090
rect 31232 6056 31236 6090
rect 31172 6022 31236 6056
rect 31172 5988 31198 6022
rect 31232 5988 31236 6022
rect 31172 5934 31236 5988
<< nsubdiff >>
rect -4792 8306 -4728 8360
rect -4792 8272 -4788 8306
rect -4754 8272 -4728 8306
rect -4792 8238 -4728 8272
rect -4792 8204 -4788 8238
rect -4754 8204 -4728 8238
rect -4792 8170 -4728 8204
rect -4792 8136 -4788 8170
rect -4754 8136 -4728 8170
rect -4792 8102 -4728 8136
rect -4792 8068 -4788 8102
rect -4754 8068 -4728 8102
rect -4792 8034 -4728 8068
rect -4792 8000 -4788 8034
rect -4754 8000 -4728 8034
rect -4792 7966 -4728 8000
rect -4792 7932 -4788 7966
rect -4754 7932 -4728 7966
rect -4792 7898 -4728 7932
rect -4792 7864 -4788 7898
rect -4754 7864 -4728 7898
rect -4792 7830 -4728 7864
rect -4792 7796 -4788 7830
rect -4754 7796 -4728 7830
rect -4792 7762 -4728 7796
rect -4792 7728 -4788 7762
rect -4754 7728 -4728 7762
rect -4792 7694 -4728 7728
rect -4792 7660 -4788 7694
rect -4754 7660 -4728 7694
rect -4792 7626 -4728 7660
rect -4792 7592 -4788 7626
rect -4754 7592 -4728 7626
rect -4792 7558 -4728 7592
rect -4792 7524 -4788 7558
rect -4754 7524 -4728 7558
rect -4792 7490 -4728 7524
rect -4792 7456 -4788 7490
rect -4754 7456 -4728 7490
rect -4792 7422 -4728 7456
rect -4792 7388 -4788 7422
rect -4754 7388 -4728 7422
rect -4792 7360 -4728 7388
rect -4410 8332 -4324 8360
rect -4410 8298 -4384 8332
rect -4350 8298 -4324 8332
rect -4410 8264 -4324 8298
rect -4410 8230 -4384 8264
rect -4350 8230 -4324 8264
rect -4410 8196 -4324 8230
rect -4410 8162 -4384 8196
rect -4350 8162 -4324 8196
rect -4410 8128 -4324 8162
rect -4410 8094 -4384 8128
rect -4350 8094 -4324 8128
rect -4410 8060 -4324 8094
rect -4410 8026 -4384 8060
rect -4350 8026 -4324 8060
rect -4410 7992 -4324 8026
rect -4410 7958 -4384 7992
rect -4350 7958 -4324 7992
rect -4410 7924 -4324 7958
rect -4410 7890 -4384 7924
rect -4350 7890 -4324 7924
rect -4410 7856 -4324 7890
rect -4410 7822 -4384 7856
rect -4350 7822 -4324 7856
rect -4410 7788 -4324 7822
rect -4410 7754 -4384 7788
rect -4350 7754 -4324 7788
rect -4410 7720 -4324 7754
rect -4410 7686 -4384 7720
rect -4350 7686 -4324 7720
rect -4410 7652 -4324 7686
rect -4410 7618 -4384 7652
rect -4350 7618 -4324 7652
rect -4410 7584 -4324 7618
rect -4410 7550 -4384 7584
rect -4350 7550 -4324 7584
rect -4410 7516 -4324 7550
rect -4410 7482 -4384 7516
rect -4350 7482 -4324 7516
rect -4410 7448 -4324 7482
rect -4410 7414 -4384 7448
rect -4350 7414 -4324 7448
rect -4410 7360 -4324 7414
rect -4006 8332 -3920 8360
rect -4006 8298 -3980 8332
rect -3946 8298 -3920 8332
rect -4006 8264 -3920 8298
rect -4006 8230 -3980 8264
rect -3946 8230 -3920 8264
rect -4006 8196 -3920 8230
rect -4006 8162 -3980 8196
rect -3946 8162 -3920 8196
rect -4006 8128 -3920 8162
rect -4006 8094 -3980 8128
rect -3946 8094 -3920 8128
rect -4006 8060 -3920 8094
rect -4006 8026 -3980 8060
rect -3946 8026 -3920 8060
rect -4006 7992 -3920 8026
rect -4006 7958 -3980 7992
rect -3946 7958 -3920 7992
rect -4006 7924 -3920 7958
rect -4006 7890 -3980 7924
rect -3946 7890 -3920 7924
rect -4006 7856 -3920 7890
rect -4006 7822 -3980 7856
rect -3946 7822 -3920 7856
rect -4006 7788 -3920 7822
rect -4006 7754 -3980 7788
rect -3946 7754 -3920 7788
rect -4006 7720 -3920 7754
rect -4006 7686 -3980 7720
rect -3946 7686 -3920 7720
rect -4006 7652 -3920 7686
rect -4006 7618 -3980 7652
rect -3946 7618 -3920 7652
rect -4006 7584 -3920 7618
rect -4006 7550 -3980 7584
rect -3946 7550 -3920 7584
rect -4006 7516 -3920 7550
rect -4006 7482 -3980 7516
rect -3946 7482 -3920 7516
rect -4006 7448 -3920 7482
rect -4006 7414 -3980 7448
rect -3946 7414 -3920 7448
rect -4006 7360 -3920 7414
rect -3602 8332 -3516 8360
rect -3602 8298 -3576 8332
rect -3542 8298 -3516 8332
rect -3602 8264 -3516 8298
rect -3602 8230 -3576 8264
rect -3542 8230 -3516 8264
rect -3602 8196 -3516 8230
rect -3602 8162 -3576 8196
rect -3542 8162 -3516 8196
rect -3602 8128 -3516 8162
rect -3602 8094 -3576 8128
rect -3542 8094 -3516 8128
rect -3602 8060 -3516 8094
rect -3602 8026 -3576 8060
rect -3542 8026 -3516 8060
rect -3602 7992 -3516 8026
rect -3602 7958 -3576 7992
rect -3542 7958 -3516 7992
rect -3602 7924 -3516 7958
rect -3602 7890 -3576 7924
rect -3542 7890 -3516 7924
rect -3602 7856 -3516 7890
rect -3602 7822 -3576 7856
rect -3542 7822 -3516 7856
rect -3602 7788 -3516 7822
rect -3602 7754 -3576 7788
rect -3542 7754 -3516 7788
rect -3602 7720 -3516 7754
rect -3602 7686 -3576 7720
rect -3542 7686 -3516 7720
rect -3602 7652 -3516 7686
rect -3602 7618 -3576 7652
rect -3542 7618 -3516 7652
rect -3602 7584 -3516 7618
rect -3602 7550 -3576 7584
rect -3542 7550 -3516 7584
rect -3602 7516 -3516 7550
rect -3602 7482 -3576 7516
rect -3542 7482 -3516 7516
rect -3602 7448 -3516 7482
rect -3602 7414 -3576 7448
rect -3542 7414 -3516 7448
rect -3602 7360 -3516 7414
rect -3198 8332 -3112 8360
rect -3198 8298 -3172 8332
rect -3138 8298 -3112 8332
rect -3198 8264 -3112 8298
rect -3198 8230 -3172 8264
rect -3138 8230 -3112 8264
rect -3198 8196 -3112 8230
rect -3198 8162 -3172 8196
rect -3138 8162 -3112 8196
rect -3198 8128 -3112 8162
rect -3198 8094 -3172 8128
rect -3138 8094 -3112 8128
rect -3198 8060 -3112 8094
rect -3198 8026 -3172 8060
rect -3138 8026 -3112 8060
rect -3198 7992 -3112 8026
rect -3198 7958 -3172 7992
rect -3138 7958 -3112 7992
rect -3198 7924 -3112 7958
rect -3198 7890 -3172 7924
rect -3138 7890 -3112 7924
rect -3198 7856 -3112 7890
rect -3198 7822 -3172 7856
rect -3138 7822 -3112 7856
rect -3198 7788 -3112 7822
rect -3198 7754 -3172 7788
rect -3138 7754 -3112 7788
rect -3198 7720 -3112 7754
rect -3198 7686 -3172 7720
rect -3138 7686 -3112 7720
rect -3198 7652 -3112 7686
rect -3198 7618 -3172 7652
rect -3138 7618 -3112 7652
rect -3198 7584 -3112 7618
rect -3198 7550 -3172 7584
rect -3138 7550 -3112 7584
rect -3198 7516 -3112 7550
rect -3198 7482 -3172 7516
rect -3138 7482 -3112 7516
rect -3198 7448 -3112 7482
rect -3198 7414 -3172 7448
rect -3138 7414 -3112 7448
rect -3198 7360 -3112 7414
rect -2794 8332 -2708 8360
rect -2794 8298 -2768 8332
rect -2734 8298 -2708 8332
rect -2794 8264 -2708 8298
rect -2794 8230 -2768 8264
rect -2734 8230 -2708 8264
rect -2794 8196 -2708 8230
rect -2794 8162 -2768 8196
rect -2734 8162 -2708 8196
rect -2794 8128 -2708 8162
rect -2794 8094 -2768 8128
rect -2734 8094 -2708 8128
rect -2794 8060 -2708 8094
rect -2794 8026 -2768 8060
rect -2734 8026 -2708 8060
rect -2794 7992 -2708 8026
rect -2794 7958 -2768 7992
rect -2734 7958 -2708 7992
rect -2794 7924 -2708 7958
rect -2794 7890 -2768 7924
rect -2734 7890 -2708 7924
rect -2794 7856 -2708 7890
rect -2794 7822 -2768 7856
rect -2734 7822 -2708 7856
rect -2794 7788 -2708 7822
rect -2794 7754 -2768 7788
rect -2734 7754 -2708 7788
rect -2794 7720 -2708 7754
rect -2794 7686 -2768 7720
rect -2734 7686 -2708 7720
rect -2794 7652 -2708 7686
rect -2794 7618 -2768 7652
rect -2734 7618 -2708 7652
rect -2794 7584 -2708 7618
rect -2794 7550 -2768 7584
rect -2734 7550 -2708 7584
rect -2794 7516 -2708 7550
rect -2794 7482 -2768 7516
rect -2734 7482 -2708 7516
rect -2794 7448 -2708 7482
rect -2794 7414 -2768 7448
rect -2734 7414 -2708 7448
rect -2794 7360 -2708 7414
rect -2390 8332 -2326 8360
rect -2390 8298 -2364 8332
rect -2330 8298 -2326 8332
rect -2390 8264 -2326 8298
rect -2390 8230 -2364 8264
rect -2330 8230 -2326 8264
rect -2390 8196 -2326 8230
rect -2390 8162 -2364 8196
rect -2330 8162 -2326 8196
rect -2390 8128 -2326 8162
rect -2390 8094 -2364 8128
rect -2330 8094 -2326 8128
rect -2390 8060 -2326 8094
rect -2390 8026 -2364 8060
rect -2330 8026 -2326 8060
rect -2390 7992 -2326 8026
rect -2390 7958 -2364 7992
rect -2330 7958 -2326 7992
rect -2390 7924 -2326 7958
rect -2390 7890 -2364 7924
rect -2330 7890 -2326 7924
rect -2390 7856 -2326 7890
rect -2390 7822 -2364 7856
rect -2330 7822 -2326 7856
rect -2390 7788 -2326 7822
rect -2390 7754 -2364 7788
rect -2330 7754 -2326 7788
rect -2390 7720 -2326 7754
rect -2390 7686 -2364 7720
rect -2330 7686 -2326 7720
rect -2390 7652 -2326 7686
rect -2390 7618 -2364 7652
rect -2330 7618 -2326 7652
rect -2390 7584 -2326 7618
rect -2390 7550 -2364 7584
rect -2330 7550 -2326 7584
rect -2390 7516 -2326 7550
rect -2390 7482 -2364 7516
rect -2330 7482 -2326 7516
rect -2390 7448 -2326 7482
rect -2390 7414 -2364 7448
rect -2330 7414 -2326 7448
rect -2390 7360 -2326 7414
rect 606 8356 670 8410
rect 606 8322 610 8356
rect 644 8322 670 8356
rect 606 8288 670 8322
rect 606 8254 610 8288
rect 644 8254 670 8288
rect 606 8220 670 8254
rect 606 8186 610 8220
rect 644 8186 670 8220
rect 606 8152 670 8186
rect 606 8118 610 8152
rect 644 8118 670 8152
rect 606 8084 670 8118
rect 606 8050 610 8084
rect 644 8050 670 8084
rect 606 8016 670 8050
rect 606 7982 610 8016
rect 644 7982 670 8016
rect 606 7948 670 7982
rect 606 7914 610 7948
rect 644 7914 670 7948
rect 606 7880 670 7914
rect 606 7846 610 7880
rect 644 7846 670 7880
rect 606 7812 670 7846
rect 606 7778 610 7812
rect 644 7778 670 7812
rect 606 7744 670 7778
rect 606 7710 610 7744
rect 644 7710 670 7744
rect 606 7676 670 7710
rect 606 7642 610 7676
rect 644 7642 670 7676
rect 606 7608 670 7642
rect 606 7574 610 7608
rect 644 7574 670 7608
rect 606 7540 670 7574
rect 606 7506 610 7540
rect 644 7506 670 7540
rect 606 7472 670 7506
rect 606 7438 610 7472
rect 644 7438 670 7472
rect 606 7410 670 7438
rect 988 8382 1074 8410
rect 988 8348 1014 8382
rect 1048 8348 1074 8382
rect 988 8314 1074 8348
rect 988 8280 1014 8314
rect 1048 8280 1074 8314
rect 988 8246 1074 8280
rect 988 8212 1014 8246
rect 1048 8212 1074 8246
rect 988 8178 1074 8212
rect 988 8144 1014 8178
rect 1048 8144 1074 8178
rect 988 8110 1074 8144
rect 988 8076 1014 8110
rect 1048 8076 1074 8110
rect 988 8042 1074 8076
rect 988 8008 1014 8042
rect 1048 8008 1074 8042
rect 988 7974 1074 8008
rect 988 7940 1014 7974
rect 1048 7940 1074 7974
rect 988 7906 1074 7940
rect 988 7872 1014 7906
rect 1048 7872 1074 7906
rect 988 7838 1074 7872
rect 988 7804 1014 7838
rect 1048 7804 1074 7838
rect 988 7770 1074 7804
rect 988 7736 1014 7770
rect 1048 7736 1074 7770
rect 988 7702 1074 7736
rect 988 7668 1014 7702
rect 1048 7668 1074 7702
rect 988 7634 1074 7668
rect 988 7600 1014 7634
rect 1048 7600 1074 7634
rect 988 7566 1074 7600
rect 988 7532 1014 7566
rect 1048 7532 1074 7566
rect 988 7498 1074 7532
rect 988 7464 1014 7498
rect 1048 7464 1074 7498
rect 988 7410 1074 7464
rect 1392 8382 1478 8410
rect 1392 8348 1418 8382
rect 1452 8348 1478 8382
rect 1392 8314 1478 8348
rect 1392 8280 1418 8314
rect 1452 8280 1478 8314
rect 1392 8246 1478 8280
rect 1392 8212 1418 8246
rect 1452 8212 1478 8246
rect 1392 8178 1478 8212
rect 1392 8144 1418 8178
rect 1452 8144 1478 8178
rect 1392 8110 1478 8144
rect 1392 8076 1418 8110
rect 1452 8076 1478 8110
rect 1392 8042 1478 8076
rect 1392 8008 1418 8042
rect 1452 8008 1478 8042
rect 1392 7974 1478 8008
rect 1392 7940 1418 7974
rect 1452 7940 1478 7974
rect 1392 7906 1478 7940
rect 1392 7872 1418 7906
rect 1452 7872 1478 7906
rect 1392 7838 1478 7872
rect 1392 7804 1418 7838
rect 1452 7804 1478 7838
rect 1392 7770 1478 7804
rect 1392 7736 1418 7770
rect 1452 7736 1478 7770
rect 1392 7702 1478 7736
rect 1392 7668 1418 7702
rect 1452 7668 1478 7702
rect 1392 7634 1478 7668
rect 1392 7600 1418 7634
rect 1452 7600 1478 7634
rect 1392 7566 1478 7600
rect 1392 7532 1418 7566
rect 1452 7532 1478 7566
rect 1392 7498 1478 7532
rect 1392 7464 1418 7498
rect 1452 7464 1478 7498
rect 1392 7410 1478 7464
rect 1796 8382 1882 8410
rect 1796 8348 1822 8382
rect 1856 8348 1882 8382
rect 1796 8314 1882 8348
rect 1796 8280 1822 8314
rect 1856 8280 1882 8314
rect 1796 8246 1882 8280
rect 1796 8212 1822 8246
rect 1856 8212 1882 8246
rect 1796 8178 1882 8212
rect 1796 8144 1822 8178
rect 1856 8144 1882 8178
rect 1796 8110 1882 8144
rect 1796 8076 1822 8110
rect 1856 8076 1882 8110
rect 1796 8042 1882 8076
rect 1796 8008 1822 8042
rect 1856 8008 1882 8042
rect 1796 7974 1882 8008
rect 1796 7940 1822 7974
rect 1856 7940 1882 7974
rect 1796 7906 1882 7940
rect 1796 7872 1822 7906
rect 1856 7872 1882 7906
rect 1796 7838 1882 7872
rect 1796 7804 1822 7838
rect 1856 7804 1882 7838
rect 1796 7770 1882 7804
rect 1796 7736 1822 7770
rect 1856 7736 1882 7770
rect 1796 7702 1882 7736
rect 1796 7668 1822 7702
rect 1856 7668 1882 7702
rect 1796 7634 1882 7668
rect 1796 7600 1822 7634
rect 1856 7600 1882 7634
rect 1796 7566 1882 7600
rect 1796 7532 1822 7566
rect 1856 7532 1882 7566
rect 1796 7498 1882 7532
rect 1796 7464 1822 7498
rect 1856 7464 1882 7498
rect 1796 7410 1882 7464
rect 2200 8382 2286 8410
rect 2200 8348 2226 8382
rect 2260 8348 2286 8382
rect 2200 8314 2286 8348
rect 2200 8280 2226 8314
rect 2260 8280 2286 8314
rect 2200 8246 2286 8280
rect 2200 8212 2226 8246
rect 2260 8212 2286 8246
rect 2200 8178 2286 8212
rect 2200 8144 2226 8178
rect 2260 8144 2286 8178
rect 2200 8110 2286 8144
rect 2200 8076 2226 8110
rect 2260 8076 2286 8110
rect 2200 8042 2286 8076
rect 2200 8008 2226 8042
rect 2260 8008 2286 8042
rect 2200 7974 2286 8008
rect 2200 7940 2226 7974
rect 2260 7940 2286 7974
rect 2200 7906 2286 7940
rect 2200 7872 2226 7906
rect 2260 7872 2286 7906
rect 2200 7838 2286 7872
rect 2200 7804 2226 7838
rect 2260 7804 2286 7838
rect 2200 7770 2286 7804
rect 2200 7736 2226 7770
rect 2260 7736 2286 7770
rect 2200 7702 2286 7736
rect 2200 7668 2226 7702
rect 2260 7668 2286 7702
rect 2200 7634 2286 7668
rect 2200 7600 2226 7634
rect 2260 7600 2286 7634
rect 2200 7566 2286 7600
rect 2200 7532 2226 7566
rect 2260 7532 2286 7566
rect 2200 7498 2286 7532
rect 2200 7464 2226 7498
rect 2260 7464 2286 7498
rect 2200 7410 2286 7464
rect 2604 8382 2690 8410
rect 2604 8348 2630 8382
rect 2664 8348 2690 8382
rect 2604 8314 2690 8348
rect 2604 8280 2630 8314
rect 2664 8280 2690 8314
rect 2604 8246 2690 8280
rect 2604 8212 2630 8246
rect 2664 8212 2690 8246
rect 2604 8178 2690 8212
rect 2604 8144 2630 8178
rect 2664 8144 2690 8178
rect 2604 8110 2690 8144
rect 2604 8076 2630 8110
rect 2664 8076 2690 8110
rect 2604 8042 2690 8076
rect 2604 8008 2630 8042
rect 2664 8008 2690 8042
rect 2604 7974 2690 8008
rect 2604 7940 2630 7974
rect 2664 7940 2690 7974
rect 2604 7906 2690 7940
rect 2604 7872 2630 7906
rect 2664 7872 2690 7906
rect 2604 7838 2690 7872
rect 2604 7804 2630 7838
rect 2664 7804 2690 7838
rect 2604 7770 2690 7804
rect 2604 7736 2630 7770
rect 2664 7736 2690 7770
rect 2604 7702 2690 7736
rect 2604 7668 2630 7702
rect 2664 7668 2690 7702
rect 2604 7634 2690 7668
rect 2604 7600 2630 7634
rect 2664 7600 2690 7634
rect 2604 7566 2690 7600
rect 2604 7532 2630 7566
rect 2664 7532 2690 7566
rect 2604 7498 2690 7532
rect 2604 7464 2630 7498
rect 2664 7464 2690 7498
rect 2604 7410 2690 7464
rect 3008 8382 3072 8410
rect 3008 8348 3034 8382
rect 3068 8348 3072 8382
rect 3008 8314 3072 8348
rect 3008 8280 3034 8314
rect 3068 8280 3072 8314
rect 3008 8246 3072 8280
rect 3008 8212 3034 8246
rect 3068 8212 3072 8246
rect 3008 8178 3072 8212
rect 3008 8144 3034 8178
rect 3068 8144 3072 8178
rect 3008 8110 3072 8144
rect 3008 8076 3034 8110
rect 3068 8076 3072 8110
rect 3008 8042 3072 8076
rect 3008 8008 3034 8042
rect 3068 8008 3072 8042
rect 3008 7974 3072 8008
rect 3008 7940 3034 7974
rect 3068 7940 3072 7974
rect 3008 7906 3072 7940
rect 3008 7872 3034 7906
rect 3068 7872 3072 7906
rect 3008 7838 3072 7872
rect 3008 7804 3034 7838
rect 3068 7804 3072 7838
rect 3008 7770 3072 7804
rect 3008 7736 3034 7770
rect 3068 7736 3072 7770
rect 3008 7702 3072 7736
rect 3008 7668 3034 7702
rect 3068 7668 3072 7702
rect 3008 7634 3072 7668
rect 3008 7600 3034 7634
rect 3068 7600 3072 7634
rect 3008 7566 3072 7600
rect 3008 7532 3034 7566
rect 3068 7532 3072 7566
rect 3008 7498 3072 7532
rect 3008 7464 3034 7498
rect 3068 7464 3072 7498
rect 3008 7410 3072 7464
rect 6976 8356 7040 8410
rect 6976 8322 6980 8356
rect 7014 8322 7040 8356
rect 6976 8288 7040 8322
rect 6976 8254 6980 8288
rect 7014 8254 7040 8288
rect 6976 8220 7040 8254
rect 6976 8186 6980 8220
rect 7014 8186 7040 8220
rect 6976 8152 7040 8186
rect 6976 8118 6980 8152
rect 7014 8118 7040 8152
rect 6976 8084 7040 8118
rect 6976 8050 6980 8084
rect 7014 8050 7040 8084
rect 6976 8016 7040 8050
rect 6976 7982 6980 8016
rect 7014 7982 7040 8016
rect 6976 7948 7040 7982
rect 6976 7914 6980 7948
rect 7014 7914 7040 7948
rect 6976 7880 7040 7914
rect 6976 7846 6980 7880
rect 7014 7846 7040 7880
rect 6976 7812 7040 7846
rect 6976 7778 6980 7812
rect 7014 7778 7040 7812
rect 6976 7744 7040 7778
rect 6976 7710 6980 7744
rect 7014 7710 7040 7744
rect 6976 7676 7040 7710
rect 6976 7642 6980 7676
rect 7014 7642 7040 7676
rect 6976 7608 7040 7642
rect 6976 7574 6980 7608
rect 7014 7574 7040 7608
rect 6976 7540 7040 7574
rect 6976 7506 6980 7540
rect 7014 7506 7040 7540
rect 6976 7472 7040 7506
rect 6976 7438 6980 7472
rect 7014 7438 7040 7472
rect 6976 7410 7040 7438
rect 7358 8382 7444 8410
rect 7358 8348 7384 8382
rect 7418 8348 7444 8382
rect 7358 8314 7444 8348
rect 7358 8280 7384 8314
rect 7418 8280 7444 8314
rect 7358 8246 7444 8280
rect 7358 8212 7384 8246
rect 7418 8212 7444 8246
rect 7358 8178 7444 8212
rect 7358 8144 7384 8178
rect 7418 8144 7444 8178
rect 7358 8110 7444 8144
rect 7358 8076 7384 8110
rect 7418 8076 7444 8110
rect 7358 8042 7444 8076
rect 7358 8008 7384 8042
rect 7418 8008 7444 8042
rect 7358 7974 7444 8008
rect 7358 7940 7384 7974
rect 7418 7940 7444 7974
rect 7358 7906 7444 7940
rect 7358 7872 7384 7906
rect 7418 7872 7444 7906
rect 7358 7838 7444 7872
rect 7358 7804 7384 7838
rect 7418 7804 7444 7838
rect 7358 7770 7444 7804
rect 7358 7736 7384 7770
rect 7418 7736 7444 7770
rect 7358 7702 7444 7736
rect 7358 7668 7384 7702
rect 7418 7668 7444 7702
rect 7358 7634 7444 7668
rect 7358 7600 7384 7634
rect 7418 7600 7444 7634
rect 7358 7566 7444 7600
rect 7358 7532 7384 7566
rect 7418 7532 7444 7566
rect 7358 7498 7444 7532
rect 7358 7464 7384 7498
rect 7418 7464 7444 7498
rect 7358 7410 7444 7464
rect 7762 8382 7848 8410
rect 7762 8348 7788 8382
rect 7822 8348 7848 8382
rect 7762 8314 7848 8348
rect 7762 8280 7788 8314
rect 7822 8280 7848 8314
rect 7762 8246 7848 8280
rect 7762 8212 7788 8246
rect 7822 8212 7848 8246
rect 7762 8178 7848 8212
rect 7762 8144 7788 8178
rect 7822 8144 7848 8178
rect 7762 8110 7848 8144
rect 7762 8076 7788 8110
rect 7822 8076 7848 8110
rect 7762 8042 7848 8076
rect 7762 8008 7788 8042
rect 7822 8008 7848 8042
rect 7762 7974 7848 8008
rect 7762 7940 7788 7974
rect 7822 7940 7848 7974
rect 7762 7906 7848 7940
rect 7762 7872 7788 7906
rect 7822 7872 7848 7906
rect 7762 7838 7848 7872
rect 7762 7804 7788 7838
rect 7822 7804 7848 7838
rect 7762 7770 7848 7804
rect 7762 7736 7788 7770
rect 7822 7736 7848 7770
rect 7762 7702 7848 7736
rect 7762 7668 7788 7702
rect 7822 7668 7848 7702
rect 7762 7634 7848 7668
rect 7762 7600 7788 7634
rect 7822 7600 7848 7634
rect 7762 7566 7848 7600
rect 7762 7532 7788 7566
rect 7822 7532 7848 7566
rect 7762 7498 7848 7532
rect 7762 7464 7788 7498
rect 7822 7464 7848 7498
rect 7762 7410 7848 7464
rect 8166 8382 8252 8410
rect 8166 8348 8192 8382
rect 8226 8348 8252 8382
rect 8166 8314 8252 8348
rect 8166 8280 8192 8314
rect 8226 8280 8252 8314
rect 8166 8246 8252 8280
rect 8166 8212 8192 8246
rect 8226 8212 8252 8246
rect 8166 8178 8252 8212
rect 8166 8144 8192 8178
rect 8226 8144 8252 8178
rect 8166 8110 8252 8144
rect 8166 8076 8192 8110
rect 8226 8076 8252 8110
rect 8166 8042 8252 8076
rect 8166 8008 8192 8042
rect 8226 8008 8252 8042
rect 8166 7974 8252 8008
rect 8166 7940 8192 7974
rect 8226 7940 8252 7974
rect 8166 7906 8252 7940
rect 8166 7872 8192 7906
rect 8226 7872 8252 7906
rect 8166 7838 8252 7872
rect 8166 7804 8192 7838
rect 8226 7804 8252 7838
rect 8166 7770 8252 7804
rect 8166 7736 8192 7770
rect 8226 7736 8252 7770
rect 8166 7702 8252 7736
rect 8166 7668 8192 7702
rect 8226 7668 8252 7702
rect 8166 7634 8252 7668
rect 8166 7600 8192 7634
rect 8226 7600 8252 7634
rect 8166 7566 8252 7600
rect 8166 7532 8192 7566
rect 8226 7532 8252 7566
rect 8166 7498 8252 7532
rect 8166 7464 8192 7498
rect 8226 7464 8252 7498
rect 8166 7410 8252 7464
rect 8570 8382 8656 8410
rect 8570 8348 8596 8382
rect 8630 8348 8656 8382
rect 8570 8314 8656 8348
rect 8570 8280 8596 8314
rect 8630 8280 8656 8314
rect 8570 8246 8656 8280
rect 8570 8212 8596 8246
rect 8630 8212 8656 8246
rect 8570 8178 8656 8212
rect 8570 8144 8596 8178
rect 8630 8144 8656 8178
rect 8570 8110 8656 8144
rect 8570 8076 8596 8110
rect 8630 8076 8656 8110
rect 8570 8042 8656 8076
rect 8570 8008 8596 8042
rect 8630 8008 8656 8042
rect 8570 7974 8656 8008
rect 8570 7940 8596 7974
rect 8630 7940 8656 7974
rect 8570 7906 8656 7940
rect 8570 7872 8596 7906
rect 8630 7872 8656 7906
rect 8570 7838 8656 7872
rect 8570 7804 8596 7838
rect 8630 7804 8656 7838
rect 8570 7770 8656 7804
rect 8570 7736 8596 7770
rect 8630 7736 8656 7770
rect 8570 7702 8656 7736
rect 8570 7668 8596 7702
rect 8630 7668 8656 7702
rect 8570 7634 8656 7668
rect 8570 7600 8596 7634
rect 8630 7600 8656 7634
rect 8570 7566 8656 7600
rect 8570 7532 8596 7566
rect 8630 7532 8656 7566
rect 8570 7498 8656 7532
rect 8570 7464 8596 7498
rect 8630 7464 8656 7498
rect 8570 7410 8656 7464
rect 8974 8382 9060 8410
rect 8974 8348 9000 8382
rect 9034 8348 9060 8382
rect 8974 8314 9060 8348
rect 8974 8280 9000 8314
rect 9034 8280 9060 8314
rect 8974 8246 9060 8280
rect 8974 8212 9000 8246
rect 9034 8212 9060 8246
rect 8974 8178 9060 8212
rect 8974 8144 9000 8178
rect 9034 8144 9060 8178
rect 8974 8110 9060 8144
rect 8974 8076 9000 8110
rect 9034 8076 9060 8110
rect 8974 8042 9060 8076
rect 8974 8008 9000 8042
rect 9034 8008 9060 8042
rect 8974 7974 9060 8008
rect 8974 7940 9000 7974
rect 9034 7940 9060 7974
rect 8974 7906 9060 7940
rect 8974 7872 9000 7906
rect 9034 7872 9060 7906
rect 8974 7838 9060 7872
rect 8974 7804 9000 7838
rect 9034 7804 9060 7838
rect 8974 7770 9060 7804
rect 8974 7736 9000 7770
rect 9034 7736 9060 7770
rect 8974 7702 9060 7736
rect 8974 7668 9000 7702
rect 9034 7668 9060 7702
rect 8974 7634 9060 7668
rect 8974 7600 9000 7634
rect 9034 7600 9060 7634
rect 8974 7566 9060 7600
rect 8974 7532 9000 7566
rect 9034 7532 9060 7566
rect 8974 7498 9060 7532
rect 8974 7464 9000 7498
rect 9034 7464 9060 7498
rect 8974 7410 9060 7464
rect 9378 8382 9442 8410
rect 9378 8348 9404 8382
rect 9438 8348 9442 8382
rect 9378 8314 9442 8348
rect 9378 8280 9404 8314
rect 9438 8280 9442 8314
rect 9378 8246 9442 8280
rect 9378 8212 9404 8246
rect 9438 8212 9442 8246
rect 9378 8178 9442 8212
rect 9378 8144 9404 8178
rect 9438 8144 9442 8178
rect 9378 8110 9442 8144
rect 9378 8076 9404 8110
rect 9438 8076 9442 8110
rect 9378 8042 9442 8076
rect 9378 8008 9404 8042
rect 9438 8008 9442 8042
rect 9378 7974 9442 8008
rect 9378 7940 9404 7974
rect 9438 7940 9442 7974
rect 9378 7906 9442 7940
rect 9378 7872 9404 7906
rect 9438 7872 9442 7906
rect 9378 7838 9442 7872
rect 9378 7804 9404 7838
rect 9438 7804 9442 7838
rect 9378 7770 9442 7804
rect 9378 7736 9404 7770
rect 9438 7736 9442 7770
rect 9378 7702 9442 7736
rect 9378 7668 9404 7702
rect 9438 7668 9442 7702
rect 9378 7634 9442 7668
rect 9378 7600 9404 7634
rect 9438 7600 9442 7634
rect 9378 7566 9442 7600
rect 9378 7532 9404 7566
rect 9438 7532 9442 7566
rect 9378 7498 9442 7532
rect 9378 7464 9404 7498
rect 9438 7464 9442 7498
rect 9378 7410 9442 7464
rect 13346 8356 13410 8410
rect 13346 8322 13350 8356
rect 13384 8322 13410 8356
rect 13346 8288 13410 8322
rect 13346 8254 13350 8288
rect 13384 8254 13410 8288
rect 13346 8220 13410 8254
rect 13346 8186 13350 8220
rect 13384 8186 13410 8220
rect 13346 8152 13410 8186
rect 13346 8118 13350 8152
rect 13384 8118 13410 8152
rect 13346 8084 13410 8118
rect 13346 8050 13350 8084
rect 13384 8050 13410 8084
rect 13346 8016 13410 8050
rect 13346 7982 13350 8016
rect 13384 7982 13410 8016
rect 13346 7948 13410 7982
rect 13346 7914 13350 7948
rect 13384 7914 13410 7948
rect 13346 7880 13410 7914
rect 13346 7846 13350 7880
rect 13384 7846 13410 7880
rect 13346 7812 13410 7846
rect 13346 7778 13350 7812
rect 13384 7778 13410 7812
rect 13346 7744 13410 7778
rect 13346 7710 13350 7744
rect 13384 7710 13410 7744
rect 13346 7676 13410 7710
rect 13346 7642 13350 7676
rect 13384 7642 13410 7676
rect 13346 7608 13410 7642
rect 13346 7574 13350 7608
rect 13384 7574 13410 7608
rect 13346 7540 13410 7574
rect 13346 7506 13350 7540
rect 13384 7506 13410 7540
rect 13346 7472 13410 7506
rect 13346 7438 13350 7472
rect 13384 7438 13410 7472
rect 13346 7410 13410 7438
rect 13728 8382 13814 8410
rect 13728 8348 13754 8382
rect 13788 8348 13814 8382
rect 13728 8314 13814 8348
rect 13728 8280 13754 8314
rect 13788 8280 13814 8314
rect 13728 8246 13814 8280
rect 13728 8212 13754 8246
rect 13788 8212 13814 8246
rect 13728 8178 13814 8212
rect 13728 8144 13754 8178
rect 13788 8144 13814 8178
rect 13728 8110 13814 8144
rect 13728 8076 13754 8110
rect 13788 8076 13814 8110
rect 13728 8042 13814 8076
rect 13728 8008 13754 8042
rect 13788 8008 13814 8042
rect 13728 7974 13814 8008
rect 13728 7940 13754 7974
rect 13788 7940 13814 7974
rect 13728 7906 13814 7940
rect 13728 7872 13754 7906
rect 13788 7872 13814 7906
rect 13728 7838 13814 7872
rect 13728 7804 13754 7838
rect 13788 7804 13814 7838
rect 13728 7770 13814 7804
rect 13728 7736 13754 7770
rect 13788 7736 13814 7770
rect 13728 7702 13814 7736
rect 13728 7668 13754 7702
rect 13788 7668 13814 7702
rect 13728 7634 13814 7668
rect 13728 7600 13754 7634
rect 13788 7600 13814 7634
rect 13728 7566 13814 7600
rect 13728 7532 13754 7566
rect 13788 7532 13814 7566
rect 13728 7498 13814 7532
rect 13728 7464 13754 7498
rect 13788 7464 13814 7498
rect 13728 7410 13814 7464
rect 14132 8382 14218 8410
rect 14132 8348 14158 8382
rect 14192 8348 14218 8382
rect 14132 8314 14218 8348
rect 14132 8280 14158 8314
rect 14192 8280 14218 8314
rect 14132 8246 14218 8280
rect 14132 8212 14158 8246
rect 14192 8212 14218 8246
rect 14132 8178 14218 8212
rect 14132 8144 14158 8178
rect 14192 8144 14218 8178
rect 14132 8110 14218 8144
rect 14132 8076 14158 8110
rect 14192 8076 14218 8110
rect 14132 8042 14218 8076
rect 14132 8008 14158 8042
rect 14192 8008 14218 8042
rect 14132 7974 14218 8008
rect 14132 7940 14158 7974
rect 14192 7940 14218 7974
rect 14132 7906 14218 7940
rect 14132 7872 14158 7906
rect 14192 7872 14218 7906
rect 14132 7838 14218 7872
rect 14132 7804 14158 7838
rect 14192 7804 14218 7838
rect 14132 7770 14218 7804
rect 14132 7736 14158 7770
rect 14192 7736 14218 7770
rect 14132 7702 14218 7736
rect 14132 7668 14158 7702
rect 14192 7668 14218 7702
rect 14132 7634 14218 7668
rect 14132 7600 14158 7634
rect 14192 7600 14218 7634
rect 14132 7566 14218 7600
rect 14132 7532 14158 7566
rect 14192 7532 14218 7566
rect 14132 7498 14218 7532
rect 14132 7464 14158 7498
rect 14192 7464 14218 7498
rect 14132 7410 14218 7464
rect 14536 8382 14622 8410
rect 14536 8348 14562 8382
rect 14596 8348 14622 8382
rect 14536 8314 14622 8348
rect 14536 8280 14562 8314
rect 14596 8280 14622 8314
rect 14536 8246 14622 8280
rect 14536 8212 14562 8246
rect 14596 8212 14622 8246
rect 14536 8178 14622 8212
rect 14536 8144 14562 8178
rect 14596 8144 14622 8178
rect 14536 8110 14622 8144
rect 14536 8076 14562 8110
rect 14596 8076 14622 8110
rect 14536 8042 14622 8076
rect 14536 8008 14562 8042
rect 14596 8008 14622 8042
rect 14536 7974 14622 8008
rect 14536 7940 14562 7974
rect 14596 7940 14622 7974
rect 14536 7906 14622 7940
rect 14536 7872 14562 7906
rect 14596 7872 14622 7906
rect 14536 7838 14622 7872
rect 14536 7804 14562 7838
rect 14596 7804 14622 7838
rect 14536 7770 14622 7804
rect 14536 7736 14562 7770
rect 14596 7736 14622 7770
rect 14536 7702 14622 7736
rect 14536 7668 14562 7702
rect 14596 7668 14622 7702
rect 14536 7634 14622 7668
rect 14536 7600 14562 7634
rect 14596 7600 14622 7634
rect 14536 7566 14622 7600
rect 14536 7532 14562 7566
rect 14596 7532 14622 7566
rect 14536 7498 14622 7532
rect 14536 7464 14562 7498
rect 14596 7464 14622 7498
rect 14536 7410 14622 7464
rect 14940 8382 15026 8410
rect 14940 8348 14966 8382
rect 15000 8348 15026 8382
rect 14940 8314 15026 8348
rect 14940 8280 14966 8314
rect 15000 8280 15026 8314
rect 14940 8246 15026 8280
rect 14940 8212 14966 8246
rect 15000 8212 15026 8246
rect 14940 8178 15026 8212
rect 14940 8144 14966 8178
rect 15000 8144 15026 8178
rect 14940 8110 15026 8144
rect 14940 8076 14966 8110
rect 15000 8076 15026 8110
rect 14940 8042 15026 8076
rect 14940 8008 14966 8042
rect 15000 8008 15026 8042
rect 14940 7974 15026 8008
rect 14940 7940 14966 7974
rect 15000 7940 15026 7974
rect 14940 7906 15026 7940
rect 14940 7872 14966 7906
rect 15000 7872 15026 7906
rect 14940 7838 15026 7872
rect 14940 7804 14966 7838
rect 15000 7804 15026 7838
rect 14940 7770 15026 7804
rect 14940 7736 14966 7770
rect 15000 7736 15026 7770
rect 14940 7702 15026 7736
rect 14940 7668 14966 7702
rect 15000 7668 15026 7702
rect 14940 7634 15026 7668
rect 14940 7600 14966 7634
rect 15000 7600 15026 7634
rect 14940 7566 15026 7600
rect 14940 7532 14966 7566
rect 15000 7532 15026 7566
rect 14940 7498 15026 7532
rect 14940 7464 14966 7498
rect 15000 7464 15026 7498
rect 14940 7410 15026 7464
rect 15344 8382 15430 8410
rect 15344 8348 15370 8382
rect 15404 8348 15430 8382
rect 15344 8314 15430 8348
rect 15344 8280 15370 8314
rect 15404 8280 15430 8314
rect 15344 8246 15430 8280
rect 15344 8212 15370 8246
rect 15404 8212 15430 8246
rect 15344 8178 15430 8212
rect 15344 8144 15370 8178
rect 15404 8144 15430 8178
rect 15344 8110 15430 8144
rect 15344 8076 15370 8110
rect 15404 8076 15430 8110
rect 15344 8042 15430 8076
rect 15344 8008 15370 8042
rect 15404 8008 15430 8042
rect 15344 7974 15430 8008
rect 15344 7940 15370 7974
rect 15404 7940 15430 7974
rect 15344 7906 15430 7940
rect 15344 7872 15370 7906
rect 15404 7872 15430 7906
rect 15344 7838 15430 7872
rect 15344 7804 15370 7838
rect 15404 7804 15430 7838
rect 15344 7770 15430 7804
rect 15344 7736 15370 7770
rect 15404 7736 15430 7770
rect 15344 7702 15430 7736
rect 15344 7668 15370 7702
rect 15404 7668 15430 7702
rect 15344 7634 15430 7668
rect 15344 7600 15370 7634
rect 15404 7600 15430 7634
rect 15344 7566 15430 7600
rect 15344 7532 15370 7566
rect 15404 7532 15430 7566
rect 15344 7498 15430 7532
rect 15344 7464 15370 7498
rect 15404 7464 15430 7498
rect 15344 7410 15430 7464
rect 15748 8382 15812 8410
rect 15748 8348 15774 8382
rect 15808 8348 15812 8382
rect 15748 8314 15812 8348
rect 15748 8280 15774 8314
rect 15808 8280 15812 8314
rect 15748 8246 15812 8280
rect 15748 8212 15774 8246
rect 15808 8212 15812 8246
rect 15748 8178 15812 8212
rect 15748 8144 15774 8178
rect 15808 8144 15812 8178
rect 15748 8110 15812 8144
rect 15748 8076 15774 8110
rect 15808 8076 15812 8110
rect 15748 8042 15812 8076
rect 15748 8008 15774 8042
rect 15808 8008 15812 8042
rect 15748 7974 15812 8008
rect 15748 7940 15774 7974
rect 15808 7940 15812 7974
rect 15748 7906 15812 7940
rect 15748 7872 15774 7906
rect 15808 7872 15812 7906
rect 15748 7838 15812 7872
rect 15748 7804 15774 7838
rect 15808 7804 15812 7838
rect 15748 7770 15812 7804
rect 15748 7736 15774 7770
rect 15808 7736 15812 7770
rect 15748 7702 15812 7736
rect 15748 7668 15774 7702
rect 15808 7668 15812 7702
rect 15748 7634 15812 7668
rect 15748 7600 15774 7634
rect 15808 7600 15812 7634
rect 15748 7566 15812 7600
rect 15748 7532 15774 7566
rect 15808 7532 15812 7566
rect 15748 7498 15812 7532
rect 15748 7464 15774 7498
rect 15808 7464 15812 7498
rect 15748 7410 15812 7464
rect 19716 8356 19780 8410
rect 19716 8322 19720 8356
rect 19754 8322 19780 8356
rect 19716 8288 19780 8322
rect 19716 8254 19720 8288
rect 19754 8254 19780 8288
rect 19716 8220 19780 8254
rect 19716 8186 19720 8220
rect 19754 8186 19780 8220
rect 19716 8152 19780 8186
rect 19716 8118 19720 8152
rect 19754 8118 19780 8152
rect 19716 8084 19780 8118
rect 19716 8050 19720 8084
rect 19754 8050 19780 8084
rect 19716 8016 19780 8050
rect 19716 7982 19720 8016
rect 19754 7982 19780 8016
rect 19716 7948 19780 7982
rect 19716 7914 19720 7948
rect 19754 7914 19780 7948
rect 19716 7880 19780 7914
rect 19716 7846 19720 7880
rect 19754 7846 19780 7880
rect 19716 7812 19780 7846
rect 19716 7778 19720 7812
rect 19754 7778 19780 7812
rect 19716 7744 19780 7778
rect 19716 7710 19720 7744
rect 19754 7710 19780 7744
rect 19716 7676 19780 7710
rect 19716 7642 19720 7676
rect 19754 7642 19780 7676
rect 19716 7608 19780 7642
rect 19716 7574 19720 7608
rect 19754 7574 19780 7608
rect 19716 7540 19780 7574
rect 19716 7506 19720 7540
rect 19754 7506 19780 7540
rect 19716 7472 19780 7506
rect 19716 7438 19720 7472
rect 19754 7438 19780 7472
rect 19716 7410 19780 7438
rect 20098 8382 20184 8410
rect 20098 8348 20124 8382
rect 20158 8348 20184 8382
rect 20098 8314 20184 8348
rect 20098 8280 20124 8314
rect 20158 8280 20184 8314
rect 20098 8246 20184 8280
rect 20098 8212 20124 8246
rect 20158 8212 20184 8246
rect 20098 8178 20184 8212
rect 20098 8144 20124 8178
rect 20158 8144 20184 8178
rect 20098 8110 20184 8144
rect 20098 8076 20124 8110
rect 20158 8076 20184 8110
rect 20098 8042 20184 8076
rect 20098 8008 20124 8042
rect 20158 8008 20184 8042
rect 20098 7974 20184 8008
rect 20098 7940 20124 7974
rect 20158 7940 20184 7974
rect 20098 7906 20184 7940
rect 20098 7872 20124 7906
rect 20158 7872 20184 7906
rect 20098 7838 20184 7872
rect 20098 7804 20124 7838
rect 20158 7804 20184 7838
rect 20098 7770 20184 7804
rect 20098 7736 20124 7770
rect 20158 7736 20184 7770
rect 20098 7702 20184 7736
rect 20098 7668 20124 7702
rect 20158 7668 20184 7702
rect 20098 7634 20184 7668
rect 20098 7600 20124 7634
rect 20158 7600 20184 7634
rect 20098 7566 20184 7600
rect 20098 7532 20124 7566
rect 20158 7532 20184 7566
rect 20098 7498 20184 7532
rect 20098 7464 20124 7498
rect 20158 7464 20184 7498
rect 20098 7410 20184 7464
rect 20502 8382 20588 8410
rect 20502 8348 20528 8382
rect 20562 8348 20588 8382
rect 20502 8314 20588 8348
rect 20502 8280 20528 8314
rect 20562 8280 20588 8314
rect 20502 8246 20588 8280
rect 20502 8212 20528 8246
rect 20562 8212 20588 8246
rect 20502 8178 20588 8212
rect 20502 8144 20528 8178
rect 20562 8144 20588 8178
rect 20502 8110 20588 8144
rect 20502 8076 20528 8110
rect 20562 8076 20588 8110
rect 20502 8042 20588 8076
rect 20502 8008 20528 8042
rect 20562 8008 20588 8042
rect 20502 7974 20588 8008
rect 20502 7940 20528 7974
rect 20562 7940 20588 7974
rect 20502 7906 20588 7940
rect 20502 7872 20528 7906
rect 20562 7872 20588 7906
rect 20502 7838 20588 7872
rect 20502 7804 20528 7838
rect 20562 7804 20588 7838
rect 20502 7770 20588 7804
rect 20502 7736 20528 7770
rect 20562 7736 20588 7770
rect 20502 7702 20588 7736
rect 20502 7668 20528 7702
rect 20562 7668 20588 7702
rect 20502 7634 20588 7668
rect 20502 7600 20528 7634
rect 20562 7600 20588 7634
rect 20502 7566 20588 7600
rect 20502 7532 20528 7566
rect 20562 7532 20588 7566
rect 20502 7498 20588 7532
rect 20502 7464 20528 7498
rect 20562 7464 20588 7498
rect 20502 7410 20588 7464
rect 20906 8382 20992 8410
rect 20906 8348 20932 8382
rect 20966 8348 20992 8382
rect 20906 8314 20992 8348
rect 20906 8280 20932 8314
rect 20966 8280 20992 8314
rect 20906 8246 20992 8280
rect 20906 8212 20932 8246
rect 20966 8212 20992 8246
rect 20906 8178 20992 8212
rect 20906 8144 20932 8178
rect 20966 8144 20992 8178
rect 20906 8110 20992 8144
rect 20906 8076 20932 8110
rect 20966 8076 20992 8110
rect 20906 8042 20992 8076
rect 20906 8008 20932 8042
rect 20966 8008 20992 8042
rect 20906 7974 20992 8008
rect 20906 7940 20932 7974
rect 20966 7940 20992 7974
rect 20906 7906 20992 7940
rect 20906 7872 20932 7906
rect 20966 7872 20992 7906
rect 20906 7838 20992 7872
rect 20906 7804 20932 7838
rect 20966 7804 20992 7838
rect 20906 7770 20992 7804
rect 20906 7736 20932 7770
rect 20966 7736 20992 7770
rect 20906 7702 20992 7736
rect 20906 7668 20932 7702
rect 20966 7668 20992 7702
rect 20906 7634 20992 7668
rect 20906 7600 20932 7634
rect 20966 7600 20992 7634
rect 20906 7566 20992 7600
rect 20906 7532 20932 7566
rect 20966 7532 20992 7566
rect 20906 7498 20992 7532
rect 20906 7464 20932 7498
rect 20966 7464 20992 7498
rect 20906 7410 20992 7464
rect 21310 8382 21396 8410
rect 21310 8348 21336 8382
rect 21370 8348 21396 8382
rect 21310 8314 21396 8348
rect 21310 8280 21336 8314
rect 21370 8280 21396 8314
rect 21310 8246 21396 8280
rect 21310 8212 21336 8246
rect 21370 8212 21396 8246
rect 21310 8178 21396 8212
rect 21310 8144 21336 8178
rect 21370 8144 21396 8178
rect 21310 8110 21396 8144
rect 21310 8076 21336 8110
rect 21370 8076 21396 8110
rect 21310 8042 21396 8076
rect 21310 8008 21336 8042
rect 21370 8008 21396 8042
rect 21310 7974 21396 8008
rect 21310 7940 21336 7974
rect 21370 7940 21396 7974
rect 21310 7906 21396 7940
rect 21310 7872 21336 7906
rect 21370 7872 21396 7906
rect 21310 7838 21396 7872
rect 21310 7804 21336 7838
rect 21370 7804 21396 7838
rect 21310 7770 21396 7804
rect 21310 7736 21336 7770
rect 21370 7736 21396 7770
rect 21310 7702 21396 7736
rect 21310 7668 21336 7702
rect 21370 7668 21396 7702
rect 21310 7634 21396 7668
rect 21310 7600 21336 7634
rect 21370 7600 21396 7634
rect 21310 7566 21396 7600
rect 21310 7532 21336 7566
rect 21370 7532 21396 7566
rect 21310 7498 21396 7532
rect 21310 7464 21336 7498
rect 21370 7464 21396 7498
rect 21310 7410 21396 7464
rect 21714 8382 21800 8410
rect 21714 8348 21740 8382
rect 21774 8348 21800 8382
rect 21714 8314 21800 8348
rect 21714 8280 21740 8314
rect 21774 8280 21800 8314
rect 21714 8246 21800 8280
rect 21714 8212 21740 8246
rect 21774 8212 21800 8246
rect 21714 8178 21800 8212
rect 21714 8144 21740 8178
rect 21774 8144 21800 8178
rect 21714 8110 21800 8144
rect 21714 8076 21740 8110
rect 21774 8076 21800 8110
rect 21714 8042 21800 8076
rect 21714 8008 21740 8042
rect 21774 8008 21800 8042
rect 21714 7974 21800 8008
rect 21714 7940 21740 7974
rect 21774 7940 21800 7974
rect 21714 7906 21800 7940
rect 21714 7872 21740 7906
rect 21774 7872 21800 7906
rect 21714 7838 21800 7872
rect 21714 7804 21740 7838
rect 21774 7804 21800 7838
rect 21714 7770 21800 7804
rect 21714 7736 21740 7770
rect 21774 7736 21800 7770
rect 21714 7702 21800 7736
rect 21714 7668 21740 7702
rect 21774 7668 21800 7702
rect 21714 7634 21800 7668
rect 21714 7600 21740 7634
rect 21774 7600 21800 7634
rect 21714 7566 21800 7600
rect 21714 7532 21740 7566
rect 21774 7532 21800 7566
rect 21714 7498 21800 7532
rect 21714 7464 21740 7498
rect 21774 7464 21800 7498
rect 21714 7410 21800 7464
rect 22118 8382 22182 8410
rect 22118 8348 22144 8382
rect 22178 8348 22182 8382
rect 22118 8314 22182 8348
rect 22118 8280 22144 8314
rect 22178 8280 22182 8314
rect 22118 8246 22182 8280
rect 22118 8212 22144 8246
rect 22178 8212 22182 8246
rect 22118 8178 22182 8212
rect 22118 8144 22144 8178
rect 22178 8144 22182 8178
rect 22118 8110 22182 8144
rect 22118 8076 22144 8110
rect 22178 8076 22182 8110
rect 22118 8042 22182 8076
rect 22118 8008 22144 8042
rect 22178 8008 22182 8042
rect 22118 7974 22182 8008
rect 22118 7940 22144 7974
rect 22178 7940 22182 7974
rect 22118 7906 22182 7940
rect 22118 7872 22144 7906
rect 22178 7872 22182 7906
rect 22118 7838 22182 7872
rect 22118 7804 22144 7838
rect 22178 7804 22182 7838
rect 22118 7770 22182 7804
rect 22118 7736 22144 7770
rect 22178 7736 22182 7770
rect 22118 7702 22182 7736
rect 22118 7668 22144 7702
rect 22178 7668 22182 7702
rect 22118 7634 22182 7668
rect 22118 7600 22144 7634
rect 22178 7600 22182 7634
rect 22118 7566 22182 7600
rect 22118 7532 22144 7566
rect 22178 7532 22182 7566
rect 22118 7498 22182 7532
rect 22118 7464 22144 7498
rect 22178 7464 22182 7498
rect 22118 7410 22182 7464
rect 28974 8356 29038 8410
rect 28974 8322 28978 8356
rect 29012 8322 29038 8356
rect 28974 8288 29038 8322
rect 28974 8254 28978 8288
rect 29012 8254 29038 8288
rect 28974 8220 29038 8254
rect 28974 8186 28978 8220
rect 29012 8186 29038 8220
rect 28974 8152 29038 8186
rect 28974 8118 28978 8152
rect 29012 8118 29038 8152
rect 28974 8084 29038 8118
rect 28974 8050 28978 8084
rect 29012 8050 29038 8084
rect 28974 8016 29038 8050
rect 28974 7982 28978 8016
rect 29012 7982 29038 8016
rect 28974 7948 29038 7982
rect 28974 7914 28978 7948
rect 29012 7914 29038 7948
rect 28974 7880 29038 7914
rect 28974 7846 28978 7880
rect 29012 7846 29038 7880
rect 28974 7812 29038 7846
rect 28974 7778 28978 7812
rect 29012 7778 29038 7812
rect 28974 7744 29038 7778
rect 28974 7710 28978 7744
rect 29012 7710 29038 7744
rect 28974 7676 29038 7710
rect 28974 7642 28978 7676
rect 29012 7642 29038 7676
rect 28974 7608 29038 7642
rect 28974 7574 28978 7608
rect 29012 7574 29038 7608
rect 28974 7540 29038 7574
rect 28974 7506 28978 7540
rect 29012 7506 29038 7540
rect 28974 7472 29038 7506
rect 28974 7438 28978 7472
rect 29012 7438 29038 7472
rect 28974 7410 29038 7438
rect 29356 8382 29442 8410
rect 29356 8348 29382 8382
rect 29416 8348 29442 8382
rect 29356 8314 29442 8348
rect 29356 8280 29382 8314
rect 29416 8280 29442 8314
rect 29356 8246 29442 8280
rect 29356 8212 29382 8246
rect 29416 8212 29442 8246
rect 29356 8178 29442 8212
rect 29356 8144 29382 8178
rect 29416 8144 29442 8178
rect 29356 8110 29442 8144
rect 29356 8076 29382 8110
rect 29416 8076 29442 8110
rect 29356 8042 29442 8076
rect 29356 8008 29382 8042
rect 29416 8008 29442 8042
rect 29356 7974 29442 8008
rect 29356 7940 29382 7974
rect 29416 7940 29442 7974
rect 29356 7906 29442 7940
rect 29356 7872 29382 7906
rect 29416 7872 29442 7906
rect 29356 7838 29442 7872
rect 29356 7804 29382 7838
rect 29416 7804 29442 7838
rect 29356 7770 29442 7804
rect 29356 7736 29382 7770
rect 29416 7736 29442 7770
rect 29356 7702 29442 7736
rect 29356 7668 29382 7702
rect 29416 7668 29442 7702
rect 29356 7634 29442 7668
rect 29356 7600 29382 7634
rect 29416 7600 29442 7634
rect 29356 7566 29442 7600
rect 29356 7532 29382 7566
rect 29416 7532 29442 7566
rect 29356 7498 29442 7532
rect 29356 7464 29382 7498
rect 29416 7464 29442 7498
rect 29356 7410 29442 7464
rect 29760 8382 29846 8410
rect 29760 8348 29786 8382
rect 29820 8348 29846 8382
rect 29760 8314 29846 8348
rect 29760 8280 29786 8314
rect 29820 8280 29846 8314
rect 29760 8246 29846 8280
rect 29760 8212 29786 8246
rect 29820 8212 29846 8246
rect 29760 8178 29846 8212
rect 29760 8144 29786 8178
rect 29820 8144 29846 8178
rect 29760 8110 29846 8144
rect 29760 8076 29786 8110
rect 29820 8076 29846 8110
rect 29760 8042 29846 8076
rect 29760 8008 29786 8042
rect 29820 8008 29846 8042
rect 29760 7974 29846 8008
rect 29760 7940 29786 7974
rect 29820 7940 29846 7974
rect 29760 7906 29846 7940
rect 29760 7872 29786 7906
rect 29820 7872 29846 7906
rect 29760 7838 29846 7872
rect 29760 7804 29786 7838
rect 29820 7804 29846 7838
rect 29760 7770 29846 7804
rect 29760 7736 29786 7770
rect 29820 7736 29846 7770
rect 29760 7702 29846 7736
rect 29760 7668 29786 7702
rect 29820 7668 29846 7702
rect 29760 7634 29846 7668
rect 29760 7600 29786 7634
rect 29820 7600 29846 7634
rect 29760 7566 29846 7600
rect 29760 7532 29786 7566
rect 29820 7532 29846 7566
rect 29760 7498 29846 7532
rect 29760 7464 29786 7498
rect 29820 7464 29846 7498
rect 29760 7410 29846 7464
rect 30164 8382 30250 8410
rect 30164 8348 30190 8382
rect 30224 8348 30250 8382
rect 30164 8314 30250 8348
rect 30164 8280 30190 8314
rect 30224 8280 30250 8314
rect 30164 8246 30250 8280
rect 30164 8212 30190 8246
rect 30224 8212 30250 8246
rect 30164 8178 30250 8212
rect 30164 8144 30190 8178
rect 30224 8144 30250 8178
rect 30164 8110 30250 8144
rect 30164 8076 30190 8110
rect 30224 8076 30250 8110
rect 30164 8042 30250 8076
rect 30164 8008 30190 8042
rect 30224 8008 30250 8042
rect 30164 7974 30250 8008
rect 30164 7940 30190 7974
rect 30224 7940 30250 7974
rect 30164 7906 30250 7940
rect 30164 7872 30190 7906
rect 30224 7872 30250 7906
rect 30164 7838 30250 7872
rect 30164 7804 30190 7838
rect 30224 7804 30250 7838
rect 30164 7770 30250 7804
rect 30164 7736 30190 7770
rect 30224 7736 30250 7770
rect 30164 7702 30250 7736
rect 30164 7668 30190 7702
rect 30224 7668 30250 7702
rect 30164 7634 30250 7668
rect 30164 7600 30190 7634
rect 30224 7600 30250 7634
rect 30164 7566 30250 7600
rect 30164 7532 30190 7566
rect 30224 7532 30250 7566
rect 30164 7498 30250 7532
rect 30164 7464 30190 7498
rect 30224 7464 30250 7498
rect 30164 7410 30250 7464
rect 30568 8382 30654 8410
rect 30568 8348 30594 8382
rect 30628 8348 30654 8382
rect 30568 8314 30654 8348
rect 30568 8280 30594 8314
rect 30628 8280 30654 8314
rect 30568 8246 30654 8280
rect 30568 8212 30594 8246
rect 30628 8212 30654 8246
rect 30568 8178 30654 8212
rect 30568 8144 30594 8178
rect 30628 8144 30654 8178
rect 30568 8110 30654 8144
rect 30568 8076 30594 8110
rect 30628 8076 30654 8110
rect 30568 8042 30654 8076
rect 30568 8008 30594 8042
rect 30628 8008 30654 8042
rect 30568 7974 30654 8008
rect 30568 7940 30594 7974
rect 30628 7940 30654 7974
rect 30568 7906 30654 7940
rect 30568 7872 30594 7906
rect 30628 7872 30654 7906
rect 30568 7838 30654 7872
rect 30568 7804 30594 7838
rect 30628 7804 30654 7838
rect 30568 7770 30654 7804
rect 30568 7736 30594 7770
rect 30628 7736 30654 7770
rect 30568 7702 30654 7736
rect 30568 7668 30594 7702
rect 30628 7668 30654 7702
rect 30568 7634 30654 7668
rect 30568 7600 30594 7634
rect 30628 7600 30654 7634
rect 30568 7566 30654 7600
rect 30568 7532 30594 7566
rect 30628 7532 30654 7566
rect 30568 7498 30654 7532
rect 30568 7464 30594 7498
rect 30628 7464 30654 7498
rect 30568 7410 30654 7464
rect 30972 8382 31058 8410
rect 30972 8348 30998 8382
rect 31032 8348 31058 8382
rect 30972 8314 31058 8348
rect 30972 8280 30998 8314
rect 31032 8280 31058 8314
rect 30972 8246 31058 8280
rect 30972 8212 30998 8246
rect 31032 8212 31058 8246
rect 30972 8178 31058 8212
rect 30972 8144 30998 8178
rect 31032 8144 31058 8178
rect 30972 8110 31058 8144
rect 30972 8076 30998 8110
rect 31032 8076 31058 8110
rect 30972 8042 31058 8076
rect 30972 8008 30998 8042
rect 31032 8008 31058 8042
rect 30972 7974 31058 8008
rect 30972 7940 30998 7974
rect 31032 7940 31058 7974
rect 30972 7906 31058 7940
rect 30972 7872 30998 7906
rect 31032 7872 31058 7906
rect 30972 7838 31058 7872
rect 30972 7804 30998 7838
rect 31032 7804 31058 7838
rect 30972 7770 31058 7804
rect 30972 7736 30998 7770
rect 31032 7736 31058 7770
rect 30972 7702 31058 7736
rect 30972 7668 30998 7702
rect 31032 7668 31058 7702
rect 30972 7634 31058 7668
rect 30972 7600 30998 7634
rect 31032 7600 31058 7634
rect 30972 7566 31058 7600
rect 30972 7532 30998 7566
rect 31032 7532 31058 7566
rect 30972 7498 31058 7532
rect 30972 7464 30998 7498
rect 31032 7464 31058 7498
rect 30972 7410 31058 7464
rect 31376 8382 31440 8410
rect 31376 8348 31402 8382
rect 31436 8348 31440 8382
rect 31376 8314 31440 8348
rect 31376 8280 31402 8314
rect 31436 8280 31440 8314
rect 31376 8246 31440 8280
rect 31376 8212 31402 8246
rect 31436 8212 31440 8246
rect 31376 8178 31440 8212
rect 31376 8144 31402 8178
rect 31436 8144 31440 8178
rect 31376 8110 31440 8144
rect 31376 8076 31402 8110
rect 31436 8076 31440 8110
rect 31376 8042 31440 8076
rect 31376 8008 31402 8042
rect 31436 8008 31440 8042
rect 31376 7974 31440 8008
rect 31376 7940 31402 7974
rect 31436 7940 31440 7974
rect 31376 7906 31440 7940
rect 31376 7872 31402 7906
rect 31436 7872 31440 7906
rect 31376 7838 31440 7872
rect 31376 7804 31402 7838
rect 31436 7804 31440 7838
rect 31376 7770 31440 7804
rect 31376 7736 31402 7770
rect 31436 7736 31440 7770
rect 31376 7702 31440 7736
rect 31376 7668 31402 7702
rect 31436 7668 31440 7702
rect 31376 7634 31440 7668
rect 31376 7600 31402 7634
rect 31436 7600 31440 7634
rect 31376 7566 31440 7600
rect 31376 7532 31402 7566
rect 31436 7532 31440 7566
rect 31376 7498 31440 7532
rect 31376 7464 31402 7498
rect 31436 7464 31440 7498
rect 31376 7410 31440 7464
<< psubdiffcont >>
rect -4584 6796 -4550 6830
rect -4584 6728 -4550 6762
rect -4584 6660 -4550 6694
rect -4584 6592 -4550 6626
rect -4584 6524 -4550 6558
rect -4584 6456 -4550 6490
rect -4584 6388 -4550 6422
rect -4584 6320 -4550 6354
rect -4584 6252 -4550 6286
rect -4584 6184 -4550 6218
rect -4584 6116 -4550 6150
rect -4584 6048 -4550 6082
rect -4584 5980 -4550 6014
rect -4584 5912 -4550 5946
rect -4248 6822 -4214 6856
rect -4248 6754 -4214 6788
rect -4248 6686 -4214 6720
rect -4248 6618 -4214 6652
rect -4248 6550 -4214 6584
rect -4248 6482 -4214 6516
rect -4248 6414 -4214 6448
rect -4248 6346 -4214 6380
rect -4248 6278 -4214 6312
rect -4248 6210 -4214 6244
rect -4248 6142 -4214 6176
rect -4248 6074 -4214 6108
rect -4248 6006 -4214 6040
rect -4248 5938 -4214 5972
rect -3912 6822 -3878 6856
rect -3912 6754 -3878 6788
rect -3912 6686 -3878 6720
rect -3912 6618 -3878 6652
rect -3912 6550 -3878 6584
rect -3912 6482 -3878 6516
rect -3912 6414 -3878 6448
rect -3912 6346 -3878 6380
rect -3912 6278 -3878 6312
rect -3912 6210 -3878 6244
rect -3912 6142 -3878 6176
rect -3912 6074 -3878 6108
rect -3912 6006 -3878 6040
rect -3912 5938 -3878 5972
rect -3576 6822 -3542 6856
rect -3576 6754 -3542 6788
rect -3576 6686 -3542 6720
rect -3576 6618 -3542 6652
rect -3576 6550 -3542 6584
rect -3576 6482 -3542 6516
rect -3576 6414 -3542 6448
rect -3576 6346 -3542 6380
rect -3576 6278 -3542 6312
rect -3576 6210 -3542 6244
rect -3576 6142 -3542 6176
rect -3576 6074 -3542 6108
rect -3576 6006 -3542 6040
rect -3576 5938 -3542 5972
rect -3240 6822 -3206 6856
rect -3240 6754 -3206 6788
rect -3240 6686 -3206 6720
rect -3240 6618 -3206 6652
rect -3240 6550 -3206 6584
rect -3240 6482 -3206 6516
rect -3240 6414 -3206 6448
rect -3240 6346 -3206 6380
rect -3240 6278 -3206 6312
rect -3240 6210 -3206 6244
rect -3240 6142 -3206 6176
rect -3240 6074 -3206 6108
rect -3240 6006 -3206 6040
rect -3240 5938 -3206 5972
rect -2904 6822 -2870 6856
rect -2904 6754 -2870 6788
rect -2904 6686 -2870 6720
rect -2904 6618 -2870 6652
rect -2904 6550 -2870 6584
rect -2904 6482 -2870 6516
rect -2904 6414 -2870 6448
rect -2904 6346 -2870 6380
rect -2904 6278 -2870 6312
rect -2904 6210 -2870 6244
rect -2904 6142 -2870 6176
rect -2904 6074 -2870 6108
rect -2904 6006 -2870 6040
rect -2904 5938 -2870 5972
rect -2568 6822 -2534 6856
rect -2568 6754 -2534 6788
rect -2568 6686 -2534 6720
rect -2568 6618 -2534 6652
rect -2568 6550 -2534 6584
rect -2568 6482 -2534 6516
rect -2568 6414 -2534 6448
rect -2568 6346 -2534 6380
rect -2568 6278 -2534 6312
rect -2568 6210 -2534 6244
rect -2568 6142 -2534 6176
rect -2568 6074 -2534 6108
rect -2568 6006 -2534 6040
rect -2568 5938 -2534 5972
rect 814 6846 848 6880
rect 814 6778 848 6812
rect 814 6710 848 6744
rect 814 6642 848 6676
rect 814 6574 848 6608
rect 814 6506 848 6540
rect 814 6438 848 6472
rect 814 6370 848 6404
rect 814 6302 848 6336
rect 814 6234 848 6268
rect 814 6166 848 6200
rect 814 6098 848 6132
rect 814 6030 848 6064
rect 814 5962 848 5996
rect 1150 6872 1184 6906
rect 1150 6804 1184 6838
rect 1150 6736 1184 6770
rect 1150 6668 1184 6702
rect 1150 6600 1184 6634
rect 1150 6532 1184 6566
rect 1150 6464 1184 6498
rect 1150 6396 1184 6430
rect 1150 6328 1184 6362
rect 1150 6260 1184 6294
rect 1150 6192 1184 6226
rect 1150 6124 1184 6158
rect 1150 6056 1184 6090
rect 1150 5988 1184 6022
rect 1486 6872 1520 6906
rect 1486 6804 1520 6838
rect 1486 6736 1520 6770
rect 1486 6668 1520 6702
rect 1486 6600 1520 6634
rect 1486 6532 1520 6566
rect 1486 6464 1520 6498
rect 1486 6396 1520 6430
rect 1486 6328 1520 6362
rect 1486 6260 1520 6294
rect 1486 6192 1520 6226
rect 1486 6124 1520 6158
rect 1486 6056 1520 6090
rect 1486 5988 1520 6022
rect 1822 6872 1856 6906
rect 1822 6804 1856 6838
rect 1822 6736 1856 6770
rect 1822 6668 1856 6702
rect 1822 6600 1856 6634
rect 1822 6532 1856 6566
rect 1822 6464 1856 6498
rect 1822 6396 1856 6430
rect 1822 6328 1856 6362
rect 1822 6260 1856 6294
rect 1822 6192 1856 6226
rect 1822 6124 1856 6158
rect 1822 6056 1856 6090
rect 1822 5988 1856 6022
rect 2158 6872 2192 6906
rect 2158 6804 2192 6838
rect 2158 6736 2192 6770
rect 2158 6668 2192 6702
rect 2158 6600 2192 6634
rect 2158 6532 2192 6566
rect 2158 6464 2192 6498
rect 2158 6396 2192 6430
rect 2158 6328 2192 6362
rect 2158 6260 2192 6294
rect 2158 6192 2192 6226
rect 2158 6124 2192 6158
rect 2158 6056 2192 6090
rect 2158 5988 2192 6022
rect 2494 6872 2528 6906
rect 2494 6804 2528 6838
rect 2494 6736 2528 6770
rect 2494 6668 2528 6702
rect 2494 6600 2528 6634
rect 2494 6532 2528 6566
rect 2494 6464 2528 6498
rect 2494 6396 2528 6430
rect 2494 6328 2528 6362
rect 2494 6260 2528 6294
rect 2494 6192 2528 6226
rect 2494 6124 2528 6158
rect 2494 6056 2528 6090
rect 2494 5988 2528 6022
rect 2830 6872 2864 6906
rect 2830 6804 2864 6838
rect 2830 6736 2864 6770
rect 2830 6668 2864 6702
rect 2830 6600 2864 6634
rect 2830 6532 2864 6566
rect 2830 6464 2864 6498
rect 2830 6396 2864 6430
rect 2830 6328 2864 6362
rect 2830 6260 2864 6294
rect 2830 6192 2864 6226
rect 2830 6124 2864 6158
rect 2830 6056 2864 6090
rect 2830 5988 2864 6022
rect 7184 6846 7218 6880
rect 7184 6778 7218 6812
rect 7184 6710 7218 6744
rect 7184 6642 7218 6676
rect 7184 6574 7218 6608
rect 7184 6506 7218 6540
rect 7184 6438 7218 6472
rect 7184 6370 7218 6404
rect 7184 6302 7218 6336
rect 7184 6234 7218 6268
rect 7184 6166 7218 6200
rect 7184 6098 7218 6132
rect 7184 6030 7218 6064
rect 7184 5962 7218 5996
rect 7520 6872 7554 6906
rect 7520 6804 7554 6838
rect 7520 6736 7554 6770
rect 7520 6668 7554 6702
rect 7520 6600 7554 6634
rect 7520 6532 7554 6566
rect 7520 6464 7554 6498
rect 7520 6396 7554 6430
rect 7520 6328 7554 6362
rect 7520 6260 7554 6294
rect 7520 6192 7554 6226
rect 7520 6124 7554 6158
rect 7520 6056 7554 6090
rect 7520 5988 7554 6022
rect 7856 6872 7890 6906
rect 7856 6804 7890 6838
rect 7856 6736 7890 6770
rect 7856 6668 7890 6702
rect 7856 6600 7890 6634
rect 7856 6532 7890 6566
rect 7856 6464 7890 6498
rect 7856 6396 7890 6430
rect 7856 6328 7890 6362
rect 7856 6260 7890 6294
rect 7856 6192 7890 6226
rect 7856 6124 7890 6158
rect 7856 6056 7890 6090
rect 7856 5988 7890 6022
rect 8192 6872 8226 6906
rect 8192 6804 8226 6838
rect 8192 6736 8226 6770
rect 8192 6668 8226 6702
rect 8192 6600 8226 6634
rect 8192 6532 8226 6566
rect 8192 6464 8226 6498
rect 8192 6396 8226 6430
rect 8192 6328 8226 6362
rect 8192 6260 8226 6294
rect 8192 6192 8226 6226
rect 8192 6124 8226 6158
rect 8192 6056 8226 6090
rect 8192 5988 8226 6022
rect 8528 6872 8562 6906
rect 8528 6804 8562 6838
rect 8528 6736 8562 6770
rect 8528 6668 8562 6702
rect 8528 6600 8562 6634
rect 8528 6532 8562 6566
rect 8528 6464 8562 6498
rect 8528 6396 8562 6430
rect 8528 6328 8562 6362
rect 8528 6260 8562 6294
rect 8528 6192 8562 6226
rect 8528 6124 8562 6158
rect 8528 6056 8562 6090
rect 8528 5988 8562 6022
rect 8864 6872 8898 6906
rect 8864 6804 8898 6838
rect 8864 6736 8898 6770
rect 8864 6668 8898 6702
rect 8864 6600 8898 6634
rect 8864 6532 8898 6566
rect 8864 6464 8898 6498
rect 8864 6396 8898 6430
rect 8864 6328 8898 6362
rect 8864 6260 8898 6294
rect 8864 6192 8898 6226
rect 8864 6124 8898 6158
rect 8864 6056 8898 6090
rect 8864 5988 8898 6022
rect 9200 6872 9234 6906
rect 9200 6804 9234 6838
rect 9200 6736 9234 6770
rect 9200 6668 9234 6702
rect 9200 6600 9234 6634
rect 9200 6532 9234 6566
rect 9200 6464 9234 6498
rect 9200 6396 9234 6430
rect 9200 6328 9234 6362
rect 9200 6260 9234 6294
rect 9200 6192 9234 6226
rect 9200 6124 9234 6158
rect 9200 6056 9234 6090
rect 9200 5988 9234 6022
rect 13554 6846 13588 6880
rect 13554 6778 13588 6812
rect 13554 6710 13588 6744
rect 13554 6642 13588 6676
rect 13554 6574 13588 6608
rect 13554 6506 13588 6540
rect 13554 6438 13588 6472
rect 13554 6370 13588 6404
rect 13554 6302 13588 6336
rect 13554 6234 13588 6268
rect 13554 6166 13588 6200
rect 13554 6098 13588 6132
rect 13554 6030 13588 6064
rect 13554 5962 13588 5996
rect 13890 6872 13924 6906
rect 13890 6804 13924 6838
rect 13890 6736 13924 6770
rect 13890 6668 13924 6702
rect 13890 6600 13924 6634
rect 13890 6532 13924 6566
rect 13890 6464 13924 6498
rect 13890 6396 13924 6430
rect 13890 6328 13924 6362
rect 13890 6260 13924 6294
rect 13890 6192 13924 6226
rect 13890 6124 13924 6158
rect 13890 6056 13924 6090
rect 13890 5988 13924 6022
rect 14226 6872 14260 6906
rect 14226 6804 14260 6838
rect 14226 6736 14260 6770
rect 14226 6668 14260 6702
rect 14226 6600 14260 6634
rect 14226 6532 14260 6566
rect 14226 6464 14260 6498
rect 14226 6396 14260 6430
rect 14226 6328 14260 6362
rect 14226 6260 14260 6294
rect 14226 6192 14260 6226
rect 14226 6124 14260 6158
rect 14226 6056 14260 6090
rect 14226 5988 14260 6022
rect 14562 6872 14596 6906
rect 14562 6804 14596 6838
rect 14562 6736 14596 6770
rect 14562 6668 14596 6702
rect 14562 6600 14596 6634
rect 14562 6532 14596 6566
rect 14562 6464 14596 6498
rect 14562 6396 14596 6430
rect 14562 6328 14596 6362
rect 14562 6260 14596 6294
rect 14562 6192 14596 6226
rect 14562 6124 14596 6158
rect 14562 6056 14596 6090
rect 14562 5988 14596 6022
rect 14898 6872 14932 6906
rect 14898 6804 14932 6838
rect 14898 6736 14932 6770
rect 14898 6668 14932 6702
rect 14898 6600 14932 6634
rect 14898 6532 14932 6566
rect 14898 6464 14932 6498
rect 14898 6396 14932 6430
rect 14898 6328 14932 6362
rect 14898 6260 14932 6294
rect 14898 6192 14932 6226
rect 14898 6124 14932 6158
rect 14898 6056 14932 6090
rect 14898 5988 14932 6022
rect 15234 6872 15268 6906
rect 15234 6804 15268 6838
rect 15234 6736 15268 6770
rect 15234 6668 15268 6702
rect 15234 6600 15268 6634
rect 15234 6532 15268 6566
rect 15234 6464 15268 6498
rect 15234 6396 15268 6430
rect 15234 6328 15268 6362
rect 15234 6260 15268 6294
rect 15234 6192 15268 6226
rect 15234 6124 15268 6158
rect 15234 6056 15268 6090
rect 15234 5988 15268 6022
rect 15570 6872 15604 6906
rect 15570 6804 15604 6838
rect 15570 6736 15604 6770
rect 15570 6668 15604 6702
rect 15570 6600 15604 6634
rect 15570 6532 15604 6566
rect 15570 6464 15604 6498
rect 15570 6396 15604 6430
rect 15570 6328 15604 6362
rect 15570 6260 15604 6294
rect 15570 6192 15604 6226
rect 15570 6124 15604 6158
rect 15570 6056 15604 6090
rect 15570 5988 15604 6022
rect 19924 6846 19958 6880
rect 19924 6778 19958 6812
rect 19924 6710 19958 6744
rect 19924 6642 19958 6676
rect 19924 6574 19958 6608
rect 19924 6506 19958 6540
rect 19924 6438 19958 6472
rect 19924 6370 19958 6404
rect 19924 6302 19958 6336
rect 19924 6234 19958 6268
rect 19924 6166 19958 6200
rect 19924 6098 19958 6132
rect 19924 6030 19958 6064
rect 19924 5962 19958 5996
rect 20260 6872 20294 6906
rect 20260 6804 20294 6838
rect 20260 6736 20294 6770
rect 20260 6668 20294 6702
rect 20260 6600 20294 6634
rect 20260 6532 20294 6566
rect 20260 6464 20294 6498
rect 20260 6396 20294 6430
rect 20260 6328 20294 6362
rect 20260 6260 20294 6294
rect 20260 6192 20294 6226
rect 20260 6124 20294 6158
rect 20260 6056 20294 6090
rect 20260 5988 20294 6022
rect 20596 6872 20630 6906
rect 20596 6804 20630 6838
rect 20596 6736 20630 6770
rect 20596 6668 20630 6702
rect 20596 6600 20630 6634
rect 20596 6532 20630 6566
rect 20596 6464 20630 6498
rect 20596 6396 20630 6430
rect 20596 6328 20630 6362
rect 20596 6260 20630 6294
rect 20596 6192 20630 6226
rect 20596 6124 20630 6158
rect 20596 6056 20630 6090
rect 20596 5988 20630 6022
rect 20932 6872 20966 6906
rect 20932 6804 20966 6838
rect 20932 6736 20966 6770
rect 20932 6668 20966 6702
rect 20932 6600 20966 6634
rect 20932 6532 20966 6566
rect 20932 6464 20966 6498
rect 20932 6396 20966 6430
rect 20932 6328 20966 6362
rect 20932 6260 20966 6294
rect 20932 6192 20966 6226
rect 20932 6124 20966 6158
rect 20932 6056 20966 6090
rect 20932 5988 20966 6022
rect 21268 6872 21302 6906
rect 21268 6804 21302 6838
rect 21268 6736 21302 6770
rect 21268 6668 21302 6702
rect 21268 6600 21302 6634
rect 21268 6532 21302 6566
rect 21268 6464 21302 6498
rect 21268 6396 21302 6430
rect 21268 6328 21302 6362
rect 21268 6260 21302 6294
rect 21268 6192 21302 6226
rect 21268 6124 21302 6158
rect 21268 6056 21302 6090
rect 21268 5988 21302 6022
rect 21604 6872 21638 6906
rect 21604 6804 21638 6838
rect 21604 6736 21638 6770
rect 21604 6668 21638 6702
rect 21604 6600 21638 6634
rect 21604 6532 21638 6566
rect 21604 6464 21638 6498
rect 21604 6396 21638 6430
rect 21604 6328 21638 6362
rect 21604 6260 21638 6294
rect 21604 6192 21638 6226
rect 21604 6124 21638 6158
rect 21604 6056 21638 6090
rect 21604 5988 21638 6022
rect 21940 6872 21974 6906
rect 21940 6804 21974 6838
rect 21940 6736 21974 6770
rect 21940 6668 21974 6702
rect 21940 6600 21974 6634
rect 21940 6532 21974 6566
rect 21940 6464 21974 6498
rect 21940 6396 21974 6430
rect 21940 6328 21974 6362
rect 21940 6260 21974 6294
rect 21940 6192 21974 6226
rect 21940 6124 21974 6158
rect 21940 6056 21974 6090
rect 21940 5988 21974 6022
rect 29182 6846 29216 6880
rect 29182 6778 29216 6812
rect 29182 6710 29216 6744
rect 29182 6642 29216 6676
rect 29182 6574 29216 6608
rect 29182 6506 29216 6540
rect 29182 6438 29216 6472
rect 29182 6370 29216 6404
rect 29182 6302 29216 6336
rect 29182 6234 29216 6268
rect 29182 6166 29216 6200
rect 29182 6098 29216 6132
rect 29182 6030 29216 6064
rect 29182 5962 29216 5996
rect 29518 6872 29552 6906
rect 29518 6804 29552 6838
rect 29518 6736 29552 6770
rect 29518 6668 29552 6702
rect 29518 6600 29552 6634
rect 29518 6532 29552 6566
rect 29518 6464 29552 6498
rect 29518 6396 29552 6430
rect 29518 6328 29552 6362
rect 29518 6260 29552 6294
rect 29518 6192 29552 6226
rect 29518 6124 29552 6158
rect 29518 6056 29552 6090
rect 29518 5988 29552 6022
rect 29854 6872 29888 6906
rect 29854 6804 29888 6838
rect 29854 6736 29888 6770
rect 29854 6668 29888 6702
rect 29854 6600 29888 6634
rect 29854 6532 29888 6566
rect 29854 6464 29888 6498
rect 29854 6396 29888 6430
rect 29854 6328 29888 6362
rect 29854 6260 29888 6294
rect 29854 6192 29888 6226
rect 29854 6124 29888 6158
rect 29854 6056 29888 6090
rect 29854 5988 29888 6022
rect 30190 6872 30224 6906
rect 30190 6804 30224 6838
rect 30190 6736 30224 6770
rect 30190 6668 30224 6702
rect 30190 6600 30224 6634
rect 30190 6532 30224 6566
rect 30190 6464 30224 6498
rect 30190 6396 30224 6430
rect 30190 6328 30224 6362
rect 30190 6260 30224 6294
rect 30190 6192 30224 6226
rect 30190 6124 30224 6158
rect 30190 6056 30224 6090
rect 30190 5988 30224 6022
rect 30526 6872 30560 6906
rect 30526 6804 30560 6838
rect 30526 6736 30560 6770
rect 30526 6668 30560 6702
rect 30526 6600 30560 6634
rect 30526 6532 30560 6566
rect 30526 6464 30560 6498
rect 30526 6396 30560 6430
rect 30526 6328 30560 6362
rect 30526 6260 30560 6294
rect 30526 6192 30560 6226
rect 30526 6124 30560 6158
rect 30526 6056 30560 6090
rect 30526 5988 30560 6022
rect 30862 6872 30896 6906
rect 30862 6804 30896 6838
rect 30862 6736 30896 6770
rect 30862 6668 30896 6702
rect 30862 6600 30896 6634
rect 30862 6532 30896 6566
rect 30862 6464 30896 6498
rect 30862 6396 30896 6430
rect 30862 6328 30896 6362
rect 30862 6260 30896 6294
rect 30862 6192 30896 6226
rect 30862 6124 30896 6158
rect 30862 6056 30896 6090
rect 30862 5988 30896 6022
rect 31198 6872 31232 6906
rect 31198 6804 31232 6838
rect 31198 6736 31232 6770
rect 31198 6668 31232 6702
rect 31198 6600 31232 6634
rect 31198 6532 31232 6566
rect 31198 6464 31232 6498
rect 31198 6396 31232 6430
rect 31198 6328 31232 6362
rect 31198 6260 31232 6294
rect 31198 6192 31232 6226
rect 31198 6124 31232 6158
rect 31198 6056 31232 6090
rect 31198 5988 31232 6022
<< nsubdiffcont >>
rect -4788 8272 -4754 8306
rect -4788 8204 -4754 8238
rect -4788 8136 -4754 8170
rect -4788 8068 -4754 8102
rect -4788 8000 -4754 8034
rect -4788 7932 -4754 7966
rect -4788 7864 -4754 7898
rect -4788 7796 -4754 7830
rect -4788 7728 -4754 7762
rect -4788 7660 -4754 7694
rect -4788 7592 -4754 7626
rect -4788 7524 -4754 7558
rect -4788 7456 -4754 7490
rect -4788 7388 -4754 7422
rect -4384 8298 -4350 8332
rect -4384 8230 -4350 8264
rect -4384 8162 -4350 8196
rect -4384 8094 -4350 8128
rect -4384 8026 -4350 8060
rect -4384 7958 -4350 7992
rect -4384 7890 -4350 7924
rect -4384 7822 -4350 7856
rect -4384 7754 -4350 7788
rect -4384 7686 -4350 7720
rect -4384 7618 -4350 7652
rect -4384 7550 -4350 7584
rect -4384 7482 -4350 7516
rect -4384 7414 -4350 7448
rect -3980 8298 -3946 8332
rect -3980 8230 -3946 8264
rect -3980 8162 -3946 8196
rect -3980 8094 -3946 8128
rect -3980 8026 -3946 8060
rect -3980 7958 -3946 7992
rect -3980 7890 -3946 7924
rect -3980 7822 -3946 7856
rect -3980 7754 -3946 7788
rect -3980 7686 -3946 7720
rect -3980 7618 -3946 7652
rect -3980 7550 -3946 7584
rect -3980 7482 -3946 7516
rect -3980 7414 -3946 7448
rect -3576 8298 -3542 8332
rect -3576 8230 -3542 8264
rect -3576 8162 -3542 8196
rect -3576 8094 -3542 8128
rect -3576 8026 -3542 8060
rect -3576 7958 -3542 7992
rect -3576 7890 -3542 7924
rect -3576 7822 -3542 7856
rect -3576 7754 -3542 7788
rect -3576 7686 -3542 7720
rect -3576 7618 -3542 7652
rect -3576 7550 -3542 7584
rect -3576 7482 -3542 7516
rect -3576 7414 -3542 7448
rect -3172 8298 -3138 8332
rect -3172 8230 -3138 8264
rect -3172 8162 -3138 8196
rect -3172 8094 -3138 8128
rect -3172 8026 -3138 8060
rect -3172 7958 -3138 7992
rect -3172 7890 -3138 7924
rect -3172 7822 -3138 7856
rect -3172 7754 -3138 7788
rect -3172 7686 -3138 7720
rect -3172 7618 -3138 7652
rect -3172 7550 -3138 7584
rect -3172 7482 -3138 7516
rect -3172 7414 -3138 7448
rect -2768 8298 -2734 8332
rect -2768 8230 -2734 8264
rect -2768 8162 -2734 8196
rect -2768 8094 -2734 8128
rect -2768 8026 -2734 8060
rect -2768 7958 -2734 7992
rect -2768 7890 -2734 7924
rect -2768 7822 -2734 7856
rect -2768 7754 -2734 7788
rect -2768 7686 -2734 7720
rect -2768 7618 -2734 7652
rect -2768 7550 -2734 7584
rect -2768 7482 -2734 7516
rect -2768 7414 -2734 7448
rect -2364 8298 -2330 8332
rect -2364 8230 -2330 8264
rect -2364 8162 -2330 8196
rect -2364 8094 -2330 8128
rect -2364 8026 -2330 8060
rect -2364 7958 -2330 7992
rect -2364 7890 -2330 7924
rect -2364 7822 -2330 7856
rect -2364 7754 -2330 7788
rect -2364 7686 -2330 7720
rect -2364 7618 -2330 7652
rect -2364 7550 -2330 7584
rect -2364 7482 -2330 7516
rect -2364 7414 -2330 7448
rect 610 8322 644 8356
rect 610 8254 644 8288
rect 610 8186 644 8220
rect 610 8118 644 8152
rect 610 8050 644 8084
rect 610 7982 644 8016
rect 610 7914 644 7948
rect 610 7846 644 7880
rect 610 7778 644 7812
rect 610 7710 644 7744
rect 610 7642 644 7676
rect 610 7574 644 7608
rect 610 7506 644 7540
rect 610 7438 644 7472
rect 1014 8348 1048 8382
rect 1014 8280 1048 8314
rect 1014 8212 1048 8246
rect 1014 8144 1048 8178
rect 1014 8076 1048 8110
rect 1014 8008 1048 8042
rect 1014 7940 1048 7974
rect 1014 7872 1048 7906
rect 1014 7804 1048 7838
rect 1014 7736 1048 7770
rect 1014 7668 1048 7702
rect 1014 7600 1048 7634
rect 1014 7532 1048 7566
rect 1014 7464 1048 7498
rect 1418 8348 1452 8382
rect 1418 8280 1452 8314
rect 1418 8212 1452 8246
rect 1418 8144 1452 8178
rect 1418 8076 1452 8110
rect 1418 8008 1452 8042
rect 1418 7940 1452 7974
rect 1418 7872 1452 7906
rect 1418 7804 1452 7838
rect 1418 7736 1452 7770
rect 1418 7668 1452 7702
rect 1418 7600 1452 7634
rect 1418 7532 1452 7566
rect 1418 7464 1452 7498
rect 1822 8348 1856 8382
rect 1822 8280 1856 8314
rect 1822 8212 1856 8246
rect 1822 8144 1856 8178
rect 1822 8076 1856 8110
rect 1822 8008 1856 8042
rect 1822 7940 1856 7974
rect 1822 7872 1856 7906
rect 1822 7804 1856 7838
rect 1822 7736 1856 7770
rect 1822 7668 1856 7702
rect 1822 7600 1856 7634
rect 1822 7532 1856 7566
rect 1822 7464 1856 7498
rect 2226 8348 2260 8382
rect 2226 8280 2260 8314
rect 2226 8212 2260 8246
rect 2226 8144 2260 8178
rect 2226 8076 2260 8110
rect 2226 8008 2260 8042
rect 2226 7940 2260 7974
rect 2226 7872 2260 7906
rect 2226 7804 2260 7838
rect 2226 7736 2260 7770
rect 2226 7668 2260 7702
rect 2226 7600 2260 7634
rect 2226 7532 2260 7566
rect 2226 7464 2260 7498
rect 2630 8348 2664 8382
rect 2630 8280 2664 8314
rect 2630 8212 2664 8246
rect 2630 8144 2664 8178
rect 2630 8076 2664 8110
rect 2630 8008 2664 8042
rect 2630 7940 2664 7974
rect 2630 7872 2664 7906
rect 2630 7804 2664 7838
rect 2630 7736 2664 7770
rect 2630 7668 2664 7702
rect 2630 7600 2664 7634
rect 2630 7532 2664 7566
rect 2630 7464 2664 7498
rect 3034 8348 3068 8382
rect 3034 8280 3068 8314
rect 3034 8212 3068 8246
rect 3034 8144 3068 8178
rect 3034 8076 3068 8110
rect 3034 8008 3068 8042
rect 3034 7940 3068 7974
rect 3034 7872 3068 7906
rect 3034 7804 3068 7838
rect 3034 7736 3068 7770
rect 3034 7668 3068 7702
rect 3034 7600 3068 7634
rect 3034 7532 3068 7566
rect 3034 7464 3068 7498
rect 6980 8322 7014 8356
rect 6980 8254 7014 8288
rect 6980 8186 7014 8220
rect 6980 8118 7014 8152
rect 6980 8050 7014 8084
rect 6980 7982 7014 8016
rect 6980 7914 7014 7948
rect 6980 7846 7014 7880
rect 6980 7778 7014 7812
rect 6980 7710 7014 7744
rect 6980 7642 7014 7676
rect 6980 7574 7014 7608
rect 6980 7506 7014 7540
rect 6980 7438 7014 7472
rect 7384 8348 7418 8382
rect 7384 8280 7418 8314
rect 7384 8212 7418 8246
rect 7384 8144 7418 8178
rect 7384 8076 7418 8110
rect 7384 8008 7418 8042
rect 7384 7940 7418 7974
rect 7384 7872 7418 7906
rect 7384 7804 7418 7838
rect 7384 7736 7418 7770
rect 7384 7668 7418 7702
rect 7384 7600 7418 7634
rect 7384 7532 7418 7566
rect 7384 7464 7418 7498
rect 7788 8348 7822 8382
rect 7788 8280 7822 8314
rect 7788 8212 7822 8246
rect 7788 8144 7822 8178
rect 7788 8076 7822 8110
rect 7788 8008 7822 8042
rect 7788 7940 7822 7974
rect 7788 7872 7822 7906
rect 7788 7804 7822 7838
rect 7788 7736 7822 7770
rect 7788 7668 7822 7702
rect 7788 7600 7822 7634
rect 7788 7532 7822 7566
rect 7788 7464 7822 7498
rect 8192 8348 8226 8382
rect 8192 8280 8226 8314
rect 8192 8212 8226 8246
rect 8192 8144 8226 8178
rect 8192 8076 8226 8110
rect 8192 8008 8226 8042
rect 8192 7940 8226 7974
rect 8192 7872 8226 7906
rect 8192 7804 8226 7838
rect 8192 7736 8226 7770
rect 8192 7668 8226 7702
rect 8192 7600 8226 7634
rect 8192 7532 8226 7566
rect 8192 7464 8226 7498
rect 8596 8348 8630 8382
rect 8596 8280 8630 8314
rect 8596 8212 8630 8246
rect 8596 8144 8630 8178
rect 8596 8076 8630 8110
rect 8596 8008 8630 8042
rect 8596 7940 8630 7974
rect 8596 7872 8630 7906
rect 8596 7804 8630 7838
rect 8596 7736 8630 7770
rect 8596 7668 8630 7702
rect 8596 7600 8630 7634
rect 8596 7532 8630 7566
rect 8596 7464 8630 7498
rect 9000 8348 9034 8382
rect 9000 8280 9034 8314
rect 9000 8212 9034 8246
rect 9000 8144 9034 8178
rect 9000 8076 9034 8110
rect 9000 8008 9034 8042
rect 9000 7940 9034 7974
rect 9000 7872 9034 7906
rect 9000 7804 9034 7838
rect 9000 7736 9034 7770
rect 9000 7668 9034 7702
rect 9000 7600 9034 7634
rect 9000 7532 9034 7566
rect 9000 7464 9034 7498
rect 9404 8348 9438 8382
rect 9404 8280 9438 8314
rect 9404 8212 9438 8246
rect 9404 8144 9438 8178
rect 9404 8076 9438 8110
rect 9404 8008 9438 8042
rect 9404 7940 9438 7974
rect 9404 7872 9438 7906
rect 9404 7804 9438 7838
rect 9404 7736 9438 7770
rect 9404 7668 9438 7702
rect 9404 7600 9438 7634
rect 9404 7532 9438 7566
rect 9404 7464 9438 7498
rect 13350 8322 13384 8356
rect 13350 8254 13384 8288
rect 13350 8186 13384 8220
rect 13350 8118 13384 8152
rect 13350 8050 13384 8084
rect 13350 7982 13384 8016
rect 13350 7914 13384 7948
rect 13350 7846 13384 7880
rect 13350 7778 13384 7812
rect 13350 7710 13384 7744
rect 13350 7642 13384 7676
rect 13350 7574 13384 7608
rect 13350 7506 13384 7540
rect 13350 7438 13384 7472
rect 13754 8348 13788 8382
rect 13754 8280 13788 8314
rect 13754 8212 13788 8246
rect 13754 8144 13788 8178
rect 13754 8076 13788 8110
rect 13754 8008 13788 8042
rect 13754 7940 13788 7974
rect 13754 7872 13788 7906
rect 13754 7804 13788 7838
rect 13754 7736 13788 7770
rect 13754 7668 13788 7702
rect 13754 7600 13788 7634
rect 13754 7532 13788 7566
rect 13754 7464 13788 7498
rect 14158 8348 14192 8382
rect 14158 8280 14192 8314
rect 14158 8212 14192 8246
rect 14158 8144 14192 8178
rect 14158 8076 14192 8110
rect 14158 8008 14192 8042
rect 14158 7940 14192 7974
rect 14158 7872 14192 7906
rect 14158 7804 14192 7838
rect 14158 7736 14192 7770
rect 14158 7668 14192 7702
rect 14158 7600 14192 7634
rect 14158 7532 14192 7566
rect 14158 7464 14192 7498
rect 14562 8348 14596 8382
rect 14562 8280 14596 8314
rect 14562 8212 14596 8246
rect 14562 8144 14596 8178
rect 14562 8076 14596 8110
rect 14562 8008 14596 8042
rect 14562 7940 14596 7974
rect 14562 7872 14596 7906
rect 14562 7804 14596 7838
rect 14562 7736 14596 7770
rect 14562 7668 14596 7702
rect 14562 7600 14596 7634
rect 14562 7532 14596 7566
rect 14562 7464 14596 7498
rect 14966 8348 15000 8382
rect 14966 8280 15000 8314
rect 14966 8212 15000 8246
rect 14966 8144 15000 8178
rect 14966 8076 15000 8110
rect 14966 8008 15000 8042
rect 14966 7940 15000 7974
rect 14966 7872 15000 7906
rect 14966 7804 15000 7838
rect 14966 7736 15000 7770
rect 14966 7668 15000 7702
rect 14966 7600 15000 7634
rect 14966 7532 15000 7566
rect 14966 7464 15000 7498
rect 15370 8348 15404 8382
rect 15370 8280 15404 8314
rect 15370 8212 15404 8246
rect 15370 8144 15404 8178
rect 15370 8076 15404 8110
rect 15370 8008 15404 8042
rect 15370 7940 15404 7974
rect 15370 7872 15404 7906
rect 15370 7804 15404 7838
rect 15370 7736 15404 7770
rect 15370 7668 15404 7702
rect 15370 7600 15404 7634
rect 15370 7532 15404 7566
rect 15370 7464 15404 7498
rect 15774 8348 15808 8382
rect 15774 8280 15808 8314
rect 15774 8212 15808 8246
rect 15774 8144 15808 8178
rect 15774 8076 15808 8110
rect 15774 8008 15808 8042
rect 15774 7940 15808 7974
rect 15774 7872 15808 7906
rect 15774 7804 15808 7838
rect 15774 7736 15808 7770
rect 15774 7668 15808 7702
rect 15774 7600 15808 7634
rect 15774 7532 15808 7566
rect 15774 7464 15808 7498
rect 19720 8322 19754 8356
rect 19720 8254 19754 8288
rect 19720 8186 19754 8220
rect 19720 8118 19754 8152
rect 19720 8050 19754 8084
rect 19720 7982 19754 8016
rect 19720 7914 19754 7948
rect 19720 7846 19754 7880
rect 19720 7778 19754 7812
rect 19720 7710 19754 7744
rect 19720 7642 19754 7676
rect 19720 7574 19754 7608
rect 19720 7506 19754 7540
rect 19720 7438 19754 7472
rect 20124 8348 20158 8382
rect 20124 8280 20158 8314
rect 20124 8212 20158 8246
rect 20124 8144 20158 8178
rect 20124 8076 20158 8110
rect 20124 8008 20158 8042
rect 20124 7940 20158 7974
rect 20124 7872 20158 7906
rect 20124 7804 20158 7838
rect 20124 7736 20158 7770
rect 20124 7668 20158 7702
rect 20124 7600 20158 7634
rect 20124 7532 20158 7566
rect 20124 7464 20158 7498
rect 20528 8348 20562 8382
rect 20528 8280 20562 8314
rect 20528 8212 20562 8246
rect 20528 8144 20562 8178
rect 20528 8076 20562 8110
rect 20528 8008 20562 8042
rect 20528 7940 20562 7974
rect 20528 7872 20562 7906
rect 20528 7804 20562 7838
rect 20528 7736 20562 7770
rect 20528 7668 20562 7702
rect 20528 7600 20562 7634
rect 20528 7532 20562 7566
rect 20528 7464 20562 7498
rect 20932 8348 20966 8382
rect 20932 8280 20966 8314
rect 20932 8212 20966 8246
rect 20932 8144 20966 8178
rect 20932 8076 20966 8110
rect 20932 8008 20966 8042
rect 20932 7940 20966 7974
rect 20932 7872 20966 7906
rect 20932 7804 20966 7838
rect 20932 7736 20966 7770
rect 20932 7668 20966 7702
rect 20932 7600 20966 7634
rect 20932 7532 20966 7566
rect 20932 7464 20966 7498
rect 21336 8348 21370 8382
rect 21336 8280 21370 8314
rect 21336 8212 21370 8246
rect 21336 8144 21370 8178
rect 21336 8076 21370 8110
rect 21336 8008 21370 8042
rect 21336 7940 21370 7974
rect 21336 7872 21370 7906
rect 21336 7804 21370 7838
rect 21336 7736 21370 7770
rect 21336 7668 21370 7702
rect 21336 7600 21370 7634
rect 21336 7532 21370 7566
rect 21336 7464 21370 7498
rect 21740 8348 21774 8382
rect 21740 8280 21774 8314
rect 21740 8212 21774 8246
rect 21740 8144 21774 8178
rect 21740 8076 21774 8110
rect 21740 8008 21774 8042
rect 21740 7940 21774 7974
rect 21740 7872 21774 7906
rect 21740 7804 21774 7838
rect 21740 7736 21774 7770
rect 21740 7668 21774 7702
rect 21740 7600 21774 7634
rect 21740 7532 21774 7566
rect 21740 7464 21774 7498
rect 22144 8348 22178 8382
rect 22144 8280 22178 8314
rect 22144 8212 22178 8246
rect 22144 8144 22178 8178
rect 22144 8076 22178 8110
rect 22144 8008 22178 8042
rect 22144 7940 22178 7974
rect 22144 7872 22178 7906
rect 22144 7804 22178 7838
rect 22144 7736 22178 7770
rect 22144 7668 22178 7702
rect 22144 7600 22178 7634
rect 22144 7532 22178 7566
rect 22144 7464 22178 7498
rect 28978 8322 29012 8356
rect 28978 8254 29012 8288
rect 28978 8186 29012 8220
rect 28978 8118 29012 8152
rect 28978 8050 29012 8084
rect 28978 7982 29012 8016
rect 28978 7914 29012 7948
rect 28978 7846 29012 7880
rect 28978 7778 29012 7812
rect 28978 7710 29012 7744
rect 28978 7642 29012 7676
rect 28978 7574 29012 7608
rect 28978 7506 29012 7540
rect 28978 7438 29012 7472
rect 29382 8348 29416 8382
rect 29382 8280 29416 8314
rect 29382 8212 29416 8246
rect 29382 8144 29416 8178
rect 29382 8076 29416 8110
rect 29382 8008 29416 8042
rect 29382 7940 29416 7974
rect 29382 7872 29416 7906
rect 29382 7804 29416 7838
rect 29382 7736 29416 7770
rect 29382 7668 29416 7702
rect 29382 7600 29416 7634
rect 29382 7532 29416 7566
rect 29382 7464 29416 7498
rect 29786 8348 29820 8382
rect 29786 8280 29820 8314
rect 29786 8212 29820 8246
rect 29786 8144 29820 8178
rect 29786 8076 29820 8110
rect 29786 8008 29820 8042
rect 29786 7940 29820 7974
rect 29786 7872 29820 7906
rect 29786 7804 29820 7838
rect 29786 7736 29820 7770
rect 29786 7668 29820 7702
rect 29786 7600 29820 7634
rect 29786 7532 29820 7566
rect 29786 7464 29820 7498
rect 30190 8348 30224 8382
rect 30190 8280 30224 8314
rect 30190 8212 30224 8246
rect 30190 8144 30224 8178
rect 30190 8076 30224 8110
rect 30190 8008 30224 8042
rect 30190 7940 30224 7974
rect 30190 7872 30224 7906
rect 30190 7804 30224 7838
rect 30190 7736 30224 7770
rect 30190 7668 30224 7702
rect 30190 7600 30224 7634
rect 30190 7532 30224 7566
rect 30190 7464 30224 7498
rect 30594 8348 30628 8382
rect 30594 8280 30628 8314
rect 30594 8212 30628 8246
rect 30594 8144 30628 8178
rect 30594 8076 30628 8110
rect 30594 8008 30628 8042
rect 30594 7940 30628 7974
rect 30594 7872 30628 7906
rect 30594 7804 30628 7838
rect 30594 7736 30628 7770
rect 30594 7668 30628 7702
rect 30594 7600 30628 7634
rect 30594 7532 30628 7566
rect 30594 7464 30628 7498
rect 30998 8348 31032 8382
rect 30998 8280 31032 8314
rect 30998 8212 31032 8246
rect 30998 8144 31032 8178
rect 30998 8076 31032 8110
rect 30998 8008 31032 8042
rect 30998 7940 31032 7974
rect 30998 7872 31032 7906
rect 30998 7804 31032 7838
rect 30998 7736 31032 7770
rect 30998 7668 31032 7702
rect 30998 7600 31032 7634
rect 30998 7532 31032 7566
rect 30998 7464 31032 7498
rect 31402 8348 31436 8382
rect 31402 8280 31436 8314
rect 31402 8212 31436 8246
rect 31402 8144 31436 8178
rect 31402 8076 31436 8110
rect 31402 8008 31436 8042
rect 31402 7940 31436 7974
rect 31402 7872 31436 7906
rect 31402 7804 31436 7838
rect 31402 7736 31436 7770
rect 31402 7668 31436 7702
rect 31402 7600 31436 7634
rect 31402 7532 31436 7566
rect 31402 7464 31436 7498
<< poly >>
rect -4668 8441 -4598 8457
rect -4668 8407 -4652 8441
rect -4614 8407 -4598 8441
rect -4668 8360 -4598 8407
rect -4540 8441 -4470 8457
rect -4540 8407 -4524 8441
rect -4486 8407 -4470 8441
rect -4540 8360 -4470 8407
rect -4264 8441 -4194 8457
rect -4264 8407 -4248 8441
rect -4210 8407 -4194 8441
rect -4264 8360 -4194 8407
rect -4136 8441 -4066 8457
rect -4136 8407 -4120 8441
rect -4082 8407 -4066 8441
rect -4136 8360 -4066 8407
rect -3860 8441 -3790 8457
rect -3860 8407 -3844 8441
rect -3806 8407 -3790 8441
rect -3860 8360 -3790 8407
rect -3732 8441 -3662 8457
rect -3732 8407 -3716 8441
rect -3678 8407 -3662 8441
rect -3732 8360 -3662 8407
rect -3456 8441 -3386 8457
rect -3456 8407 -3440 8441
rect -3402 8407 -3386 8441
rect -3456 8360 -3386 8407
rect -3328 8441 -3258 8457
rect -3328 8407 -3312 8441
rect -3274 8407 -3258 8441
rect -3328 8360 -3258 8407
rect -3052 8441 -2982 8457
rect -3052 8407 -3036 8441
rect -2998 8407 -2982 8441
rect -3052 8360 -2982 8407
rect -2924 8441 -2854 8457
rect -2924 8407 -2908 8441
rect -2870 8407 -2854 8441
rect -2924 8360 -2854 8407
rect -2648 8441 -2578 8457
rect -2648 8407 -2632 8441
rect -2594 8407 -2578 8441
rect -2648 8360 -2578 8407
rect -2520 8441 -2450 8457
rect -2520 8407 -2504 8441
rect -2466 8407 -2450 8441
rect 730 8410 800 8436
rect 858 8410 928 8436
rect 1134 8410 1204 8436
rect 1262 8410 1332 8436
rect 1538 8410 1608 8436
rect 1666 8410 1736 8436
rect 1942 8410 2012 8436
rect 2070 8410 2140 8436
rect 2346 8410 2416 8436
rect 2474 8410 2544 8436
rect 2750 8410 2820 8436
rect 2878 8410 2948 8436
rect 7100 8410 7170 8436
rect 7228 8410 7298 8436
rect 7504 8410 7574 8436
rect 7632 8410 7702 8436
rect 7908 8410 7978 8436
rect 8036 8410 8106 8436
rect 8312 8410 8382 8436
rect 8440 8410 8510 8436
rect 8716 8410 8786 8436
rect 8844 8410 8914 8436
rect 9120 8410 9190 8436
rect 9248 8410 9318 8436
rect 13470 8410 13540 8436
rect 13598 8410 13668 8436
rect 13874 8410 13944 8436
rect 14002 8410 14072 8436
rect 14278 8410 14348 8436
rect 14406 8410 14476 8436
rect 14682 8410 14752 8436
rect 14810 8410 14880 8436
rect 15086 8410 15156 8436
rect 15214 8410 15284 8436
rect 15490 8410 15560 8436
rect 15618 8410 15688 8436
rect 19840 8410 19910 8436
rect 19968 8410 20038 8436
rect 20244 8410 20314 8436
rect 20372 8410 20442 8436
rect 20648 8410 20718 8436
rect 20776 8410 20846 8436
rect 21052 8410 21122 8436
rect 21180 8410 21250 8436
rect 21456 8410 21526 8436
rect 21584 8410 21654 8436
rect 21860 8410 21930 8436
rect 21988 8410 22058 8436
rect 29098 8410 29168 8436
rect 29226 8410 29296 8436
rect 29502 8410 29572 8436
rect 29630 8410 29700 8436
rect 29906 8410 29976 8436
rect 30034 8410 30104 8436
rect 30310 8410 30380 8436
rect 30438 8410 30508 8436
rect 30714 8410 30784 8436
rect 30842 8410 30912 8436
rect 31118 8410 31188 8436
rect 31246 8410 31316 8436
rect -2520 8360 -2450 8407
rect 730 7363 800 7410
rect -4668 7313 -4598 7360
rect -4668 7279 -4652 7313
rect -4614 7279 -4598 7313
rect -4668 7263 -4598 7279
rect -4540 7313 -4470 7360
rect -4540 7279 -4524 7313
rect -4486 7279 -4470 7313
rect -4540 7263 -4470 7279
rect -4264 7313 -4194 7360
rect -4264 7279 -4248 7313
rect -4210 7279 -4194 7313
rect -4264 7263 -4194 7279
rect -4136 7313 -4066 7360
rect -4136 7279 -4120 7313
rect -4082 7279 -4066 7313
rect -4136 7263 -4066 7279
rect -3860 7313 -3790 7360
rect -3860 7279 -3844 7313
rect -3806 7279 -3790 7313
rect -3860 7263 -3790 7279
rect -3732 7313 -3662 7360
rect -3732 7279 -3716 7313
rect -3678 7279 -3662 7313
rect -3732 7263 -3662 7279
rect -3456 7313 -3386 7360
rect -3456 7279 -3440 7313
rect -3402 7279 -3386 7313
rect -3456 7263 -3386 7279
rect -3328 7313 -3258 7360
rect -3328 7279 -3312 7313
rect -3274 7279 -3258 7313
rect -3328 7263 -3258 7279
rect -3052 7313 -2982 7360
rect -3052 7279 -3036 7313
rect -2998 7279 -2982 7313
rect -3052 7263 -2982 7279
rect -2924 7313 -2854 7360
rect -2924 7279 -2908 7313
rect -2870 7279 -2854 7313
rect -2924 7263 -2854 7279
rect -2648 7313 -2578 7360
rect -2648 7279 -2632 7313
rect -2594 7279 -2578 7313
rect -2648 7263 -2578 7279
rect -2520 7313 -2450 7360
rect 730 7329 746 7363
rect 784 7329 800 7363
rect 730 7313 800 7329
rect 858 7363 928 7410
rect 858 7329 874 7363
rect 912 7329 928 7363
rect 858 7313 928 7329
rect 1134 7363 1204 7410
rect 1134 7329 1150 7363
rect 1188 7329 1204 7363
rect 1134 7313 1204 7329
rect 1262 7363 1332 7410
rect 1262 7329 1278 7363
rect 1316 7329 1332 7363
rect 1262 7313 1332 7329
rect 1538 7363 1608 7410
rect 1538 7329 1554 7363
rect 1592 7329 1608 7363
rect 1538 7313 1608 7329
rect 1666 7363 1736 7410
rect 1666 7329 1682 7363
rect 1720 7329 1736 7363
rect 1666 7313 1736 7329
rect 1942 7363 2012 7410
rect 1942 7329 1958 7363
rect 1996 7329 2012 7363
rect 1942 7313 2012 7329
rect 2070 7363 2140 7410
rect 2070 7329 2086 7363
rect 2124 7329 2140 7363
rect 2070 7313 2140 7329
rect 2346 7363 2416 7410
rect 2346 7329 2362 7363
rect 2400 7329 2416 7363
rect 2346 7313 2416 7329
rect 2474 7363 2544 7410
rect 2474 7329 2490 7363
rect 2528 7329 2544 7363
rect 2474 7313 2544 7329
rect 2750 7363 2820 7410
rect 2750 7329 2766 7363
rect 2804 7329 2820 7363
rect 2750 7313 2820 7329
rect 2878 7363 2948 7410
rect 2878 7329 2894 7363
rect 2932 7329 2948 7363
rect 2878 7313 2948 7329
rect 7100 7363 7170 7410
rect 7100 7329 7116 7363
rect 7154 7329 7170 7363
rect 7100 7313 7170 7329
rect 7228 7363 7298 7410
rect 7228 7329 7244 7363
rect 7282 7329 7298 7363
rect 7228 7313 7298 7329
rect 7504 7363 7574 7410
rect 7504 7329 7520 7363
rect 7558 7329 7574 7363
rect 7504 7313 7574 7329
rect 7632 7363 7702 7410
rect 7632 7329 7648 7363
rect 7686 7329 7702 7363
rect 7632 7313 7702 7329
rect 7908 7363 7978 7410
rect 7908 7329 7924 7363
rect 7962 7329 7978 7363
rect 7908 7313 7978 7329
rect 8036 7363 8106 7410
rect 8036 7329 8052 7363
rect 8090 7329 8106 7363
rect 8036 7313 8106 7329
rect 8312 7363 8382 7410
rect 8312 7329 8328 7363
rect 8366 7329 8382 7363
rect 8312 7313 8382 7329
rect 8440 7363 8510 7410
rect 8440 7329 8456 7363
rect 8494 7329 8510 7363
rect 8440 7313 8510 7329
rect 8716 7363 8786 7410
rect 8716 7329 8732 7363
rect 8770 7329 8786 7363
rect 8716 7313 8786 7329
rect 8844 7363 8914 7410
rect 8844 7329 8860 7363
rect 8898 7329 8914 7363
rect 8844 7313 8914 7329
rect 9120 7363 9190 7410
rect 9120 7329 9136 7363
rect 9174 7329 9190 7363
rect 9120 7313 9190 7329
rect 9248 7363 9318 7410
rect 9248 7329 9264 7363
rect 9302 7329 9318 7363
rect 9248 7313 9318 7329
rect 13470 7363 13540 7410
rect 13470 7329 13486 7363
rect 13524 7329 13540 7363
rect 13470 7313 13540 7329
rect 13598 7363 13668 7410
rect 13598 7329 13614 7363
rect 13652 7329 13668 7363
rect 13598 7313 13668 7329
rect 13874 7363 13944 7410
rect 13874 7329 13890 7363
rect 13928 7329 13944 7363
rect 13874 7313 13944 7329
rect 14002 7363 14072 7410
rect 14002 7329 14018 7363
rect 14056 7329 14072 7363
rect 14002 7313 14072 7329
rect 14278 7363 14348 7410
rect 14278 7329 14294 7363
rect 14332 7329 14348 7363
rect 14278 7313 14348 7329
rect 14406 7363 14476 7410
rect 14406 7329 14422 7363
rect 14460 7329 14476 7363
rect 14406 7313 14476 7329
rect 14682 7363 14752 7410
rect 14682 7329 14698 7363
rect 14736 7329 14752 7363
rect 14682 7313 14752 7329
rect 14810 7363 14880 7410
rect 14810 7329 14826 7363
rect 14864 7329 14880 7363
rect 14810 7313 14880 7329
rect 15086 7363 15156 7410
rect 15086 7329 15102 7363
rect 15140 7329 15156 7363
rect 15086 7313 15156 7329
rect 15214 7363 15284 7410
rect 15214 7329 15230 7363
rect 15268 7329 15284 7363
rect 15214 7313 15284 7329
rect 15490 7363 15560 7410
rect 15490 7329 15506 7363
rect 15544 7329 15560 7363
rect 15490 7313 15560 7329
rect 15618 7363 15688 7410
rect 15618 7329 15634 7363
rect 15672 7329 15688 7363
rect 15618 7313 15688 7329
rect 19840 7363 19910 7410
rect 19840 7329 19856 7363
rect 19894 7329 19910 7363
rect 19840 7313 19910 7329
rect 19968 7363 20038 7410
rect 19968 7329 19984 7363
rect 20022 7329 20038 7363
rect 19968 7313 20038 7329
rect 20244 7363 20314 7410
rect 20244 7329 20260 7363
rect 20298 7329 20314 7363
rect 20244 7313 20314 7329
rect 20372 7363 20442 7410
rect 20372 7329 20388 7363
rect 20426 7329 20442 7363
rect 20372 7313 20442 7329
rect 20648 7363 20718 7410
rect 20648 7329 20664 7363
rect 20702 7329 20718 7363
rect 20648 7313 20718 7329
rect 20776 7363 20846 7410
rect 20776 7329 20792 7363
rect 20830 7329 20846 7363
rect 20776 7313 20846 7329
rect 21052 7363 21122 7410
rect 21052 7329 21068 7363
rect 21106 7329 21122 7363
rect 21052 7313 21122 7329
rect 21180 7363 21250 7410
rect 21180 7329 21196 7363
rect 21234 7329 21250 7363
rect 21180 7313 21250 7329
rect 21456 7363 21526 7410
rect 21456 7329 21472 7363
rect 21510 7329 21526 7363
rect 21456 7313 21526 7329
rect 21584 7363 21654 7410
rect 21584 7329 21600 7363
rect 21638 7329 21654 7363
rect 21584 7313 21654 7329
rect 21860 7363 21930 7410
rect 21860 7329 21876 7363
rect 21914 7329 21930 7363
rect 21860 7313 21930 7329
rect 21988 7363 22058 7410
rect 21988 7329 22004 7363
rect 22042 7329 22058 7363
rect 21988 7313 22058 7329
rect 29098 7363 29168 7410
rect 29098 7329 29114 7363
rect 29152 7329 29168 7363
rect 29098 7313 29168 7329
rect 29226 7363 29296 7410
rect 29226 7329 29242 7363
rect 29280 7329 29296 7363
rect 29226 7313 29296 7329
rect 29502 7363 29572 7410
rect 29502 7329 29518 7363
rect 29556 7329 29572 7363
rect 29502 7313 29572 7329
rect 29630 7363 29700 7410
rect 29630 7329 29646 7363
rect 29684 7329 29700 7363
rect 29630 7313 29700 7329
rect 29906 7363 29976 7410
rect 29906 7329 29922 7363
rect 29960 7329 29976 7363
rect 29906 7313 29976 7329
rect 30034 7363 30104 7410
rect 30034 7329 30050 7363
rect 30088 7329 30104 7363
rect 30034 7313 30104 7329
rect 30310 7363 30380 7410
rect 30310 7329 30326 7363
rect 30364 7329 30380 7363
rect 30310 7313 30380 7329
rect 30438 7363 30508 7410
rect 30438 7329 30454 7363
rect 30492 7329 30508 7363
rect 30438 7313 30508 7329
rect 30714 7363 30784 7410
rect 30714 7329 30730 7363
rect 30768 7329 30784 7363
rect 30714 7313 30784 7329
rect 30842 7363 30912 7410
rect 30842 7329 30858 7363
rect 30896 7329 30912 7363
rect 30842 7313 30912 7329
rect 31118 7363 31188 7410
rect 31118 7329 31134 7363
rect 31172 7329 31188 7363
rect 31118 7313 31188 7329
rect 31246 7363 31316 7410
rect 31246 7329 31262 7363
rect 31300 7329 31316 7363
rect 31246 7313 31316 7329
rect -2520 7279 -2504 7313
rect -2466 7279 -2450 7313
rect -2520 7263 -2450 7279
rect 919 7006 1079 7022
rect 919 6972 935 7006
rect 969 6972 1029 7006
rect 1063 6972 1079 7006
rect -4479 6956 -4319 6972
rect -4479 6922 -4463 6956
rect -4429 6922 -4369 6956
rect -4335 6922 -4319 6956
rect -4479 6906 -4319 6922
rect -4143 6956 -3983 6972
rect -4143 6922 -4127 6956
rect -4093 6922 -4033 6956
rect -3999 6922 -3983 6956
rect -4143 6906 -3983 6922
rect -3807 6956 -3647 6972
rect -3807 6922 -3791 6956
rect -3757 6922 -3697 6956
rect -3663 6922 -3647 6956
rect -3807 6906 -3647 6922
rect -3471 6956 -3311 6972
rect -3471 6922 -3455 6956
rect -3421 6922 -3361 6956
rect -3327 6922 -3311 6956
rect -3471 6906 -3311 6922
rect -3135 6956 -2975 6972
rect -3135 6922 -3119 6956
rect -3085 6922 -3025 6956
rect -2991 6922 -2975 6956
rect -3135 6906 -2975 6922
rect -2799 6956 -2639 6972
rect 919 6956 1079 6972
rect 1255 7006 1415 7022
rect 1255 6972 1271 7006
rect 1305 6972 1365 7006
rect 1399 6972 1415 7006
rect 1255 6956 1415 6972
rect 1591 7006 1751 7022
rect 1591 6972 1607 7006
rect 1641 6972 1701 7006
rect 1735 6972 1751 7006
rect 1591 6956 1751 6972
rect 1927 7006 2087 7022
rect 1927 6972 1943 7006
rect 1977 6972 2037 7006
rect 2071 6972 2087 7006
rect 1927 6956 2087 6972
rect 2263 7006 2423 7022
rect 2263 6972 2279 7006
rect 2313 6972 2373 7006
rect 2407 6972 2423 7006
rect 2263 6956 2423 6972
rect 2599 7006 2759 7022
rect 2599 6972 2615 7006
rect 2649 6972 2709 7006
rect 2743 6972 2759 7006
rect 2599 6956 2759 6972
rect 7289 7006 7449 7022
rect 7289 6972 7305 7006
rect 7339 6972 7399 7006
rect 7433 6972 7449 7006
rect 7289 6956 7449 6972
rect 7625 7006 7785 7022
rect 7625 6972 7641 7006
rect 7675 6972 7735 7006
rect 7769 6972 7785 7006
rect 7625 6956 7785 6972
rect 7961 7006 8121 7022
rect 7961 6972 7977 7006
rect 8011 6972 8071 7006
rect 8105 6972 8121 7006
rect 7961 6956 8121 6972
rect 8297 7006 8457 7022
rect 8297 6972 8313 7006
rect 8347 6972 8407 7006
rect 8441 6972 8457 7006
rect 8297 6956 8457 6972
rect 8633 7006 8793 7022
rect 8633 6972 8649 7006
rect 8683 6972 8743 7006
rect 8777 6972 8793 7006
rect 8633 6956 8793 6972
rect 8969 7006 9129 7022
rect 8969 6972 8985 7006
rect 9019 6972 9079 7006
rect 9113 6972 9129 7006
rect 8969 6956 9129 6972
rect 13659 7006 13819 7022
rect 13659 6972 13675 7006
rect 13709 6972 13769 7006
rect 13803 6972 13819 7006
rect 13659 6956 13819 6972
rect 13995 7006 14155 7022
rect 13995 6972 14011 7006
rect 14045 6972 14105 7006
rect 14139 6972 14155 7006
rect 13995 6956 14155 6972
rect 14331 7006 14491 7022
rect 14331 6972 14347 7006
rect 14381 6972 14441 7006
rect 14475 6972 14491 7006
rect 14331 6956 14491 6972
rect 14667 7006 14827 7022
rect 14667 6972 14683 7006
rect 14717 6972 14777 7006
rect 14811 6972 14827 7006
rect 14667 6956 14827 6972
rect 15003 7006 15163 7022
rect 15003 6972 15019 7006
rect 15053 6972 15113 7006
rect 15147 6972 15163 7006
rect 15003 6956 15163 6972
rect 15339 7006 15499 7022
rect 15339 6972 15355 7006
rect 15389 6972 15449 7006
rect 15483 6972 15499 7006
rect 15339 6956 15499 6972
rect 20029 7006 20189 7022
rect 20029 6972 20045 7006
rect 20079 6972 20139 7006
rect 20173 6972 20189 7006
rect 20029 6956 20189 6972
rect 20365 7006 20525 7022
rect 20365 6972 20381 7006
rect 20415 6972 20475 7006
rect 20509 6972 20525 7006
rect 20365 6956 20525 6972
rect 20701 7006 20861 7022
rect 20701 6972 20717 7006
rect 20751 6972 20811 7006
rect 20845 6972 20861 7006
rect 20701 6956 20861 6972
rect 21037 7006 21197 7022
rect 21037 6972 21053 7006
rect 21087 6972 21147 7006
rect 21181 6972 21197 7006
rect 21037 6956 21197 6972
rect 21373 7006 21533 7022
rect 21373 6972 21389 7006
rect 21423 6972 21483 7006
rect 21517 6972 21533 7006
rect 21373 6956 21533 6972
rect 21709 7006 21869 7022
rect 21709 6972 21725 7006
rect 21759 6972 21819 7006
rect 21853 6972 21869 7006
rect 21709 6956 21869 6972
rect 29287 7006 29447 7022
rect 29287 6972 29303 7006
rect 29337 6972 29397 7006
rect 29431 6972 29447 7006
rect 29287 6956 29447 6972
rect 29623 7006 29783 7022
rect 29623 6972 29639 7006
rect 29673 6972 29733 7006
rect 29767 6972 29783 7006
rect 29623 6956 29783 6972
rect 29959 7006 30119 7022
rect 29959 6972 29975 7006
rect 30009 6972 30069 7006
rect 30103 6972 30119 7006
rect 29959 6956 30119 6972
rect 30295 7006 30455 7022
rect 30295 6972 30311 7006
rect 30345 6972 30405 7006
rect 30439 6972 30455 7006
rect 30295 6956 30455 6972
rect 30631 7006 30791 7022
rect 30631 6972 30647 7006
rect 30681 6972 30741 7006
rect 30775 6972 30791 7006
rect 30631 6956 30791 6972
rect 30967 7006 31127 7022
rect 30967 6972 30983 7006
rect 31017 6972 31077 7006
rect 31111 6972 31127 7006
rect 30967 6956 31127 6972
rect -2799 6922 -2783 6956
rect -2749 6922 -2689 6956
rect -2655 6922 -2639 6956
rect 934 6934 970 6956
rect 1028 6934 1064 6956
rect 1270 6934 1306 6956
rect 1364 6934 1400 6956
rect 1606 6934 1642 6956
rect 1700 6934 1736 6956
rect 1942 6934 1978 6956
rect 2036 6934 2072 6956
rect 2278 6934 2314 6956
rect 2372 6934 2408 6956
rect 2614 6934 2650 6956
rect 2708 6934 2744 6956
rect 7304 6934 7340 6956
rect 7398 6934 7434 6956
rect 7640 6934 7676 6956
rect 7734 6934 7770 6956
rect 7976 6934 8012 6956
rect 8070 6934 8106 6956
rect 8312 6934 8348 6956
rect 8406 6934 8442 6956
rect 8648 6934 8684 6956
rect 8742 6934 8778 6956
rect 8984 6934 9020 6956
rect 9078 6934 9114 6956
rect 13674 6934 13710 6956
rect 13768 6934 13804 6956
rect 14010 6934 14046 6956
rect 14104 6934 14140 6956
rect 14346 6934 14382 6956
rect 14440 6934 14476 6956
rect 14682 6934 14718 6956
rect 14776 6934 14812 6956
rect 15018 6934 15054 6956
rect 15112 6934 15148 6956
rect 15354 6934 15390 6956
rect 15448 6934 15484 6956
rect 20044 6934 20080 6956
rect 20138 6934 20174 6956
rect 20380 6934 20416 6956
rect 20474 6934 20510 6956
rect 20716 6934 20752 6956
rect 20810 6934 20846 6956
rect 21052 6934 21088 6956
rect 21146 6934 21182 6956
rect 21388 6934 21424 6956
rect 21482 6934 21518 6956
rect 21724 6934 21760 6956
rect 21818 6934 21854 6956
rect 29302 6934 29338 6956
rect 29396 6934 29432 6956
rect 29638 6934 29674 6956
rect 29732 6934 29768 6956
rect 29974 6934 30010 6956
rect 30068 6934 30104 6956
rect 30310 6934 30346 6956
rect 30404 6934 30440 6956
rect 30646 6934 30682 6956
rect 30740 6934 30776 6956
rect 30982 6934 31018 6956
rect 31076 6934 31112 6956
rect -2799 6906 -2639 6922
rect -4464 6884 -4428 6906
rect -4370 6884 -4334 6906
rect -4128 6884 -4092 6906
rect -4034 6884 -3998 6906
rect -3792 6884 -3756 6906
rect -3698 6884 -3662 6906
rect -3456 6884 -3420 6906
rect -3362 6884 -3326 6906
rect -3120 6884 -3084 6906
rect -3026 6884 -2990 6906
rect -2784 6884 -2748 6906
rect -2690 6884 -2654 6906
rect 934 5908 970 5934
rect 1028 5908 1064 5934
rect 1270 5908 1306 5934
rect 1364 5908 1400 5934
rect 1606 5908 1642 5934
rect 1700 5908 1736 5934
rect 1942 5908 1978 5934
rect 2036 5908 2072 5934
rect 2278 5908 2314 5934
rect 2372 5908 2408 5934
rect 2614 5908 2650 5934
rect 2708 5908 2744 5934
rect 7304 5908 7340 5934
rect 7398 5908 7434 5934
rect 7640 5908 7676 5934
rect 7734 5908 7770 5934
rect 7976 5908 8012 5934
rect 8070 5908 8106 5934
rect 8312 5908 8348 5934
rect 8406 5908 8442 5934
rect 8648 5908 8684 5934
rect 8742 5908 8778 5934
rect 8984 5908 9020 5934
rect 9078 5908 9114 5934
rect 13674 5908 13710 5934
rect 13768 5908 13804 5934
rect 14010 5908 14046 5934
rect 14104 5908 14140 5934
rect 14346 5908 14382 5934
rect 14440 5908 14476 5934
rect 14682 5908 14718 5934
rect 14776 5908 14812 5934
rect 15018 5908 15054 5934
rect 15112 5908 15148 5934
rect 15354 5908 15390 5934
rect 15448 5908 15484 5934
rect 20044 5908 20080 5934
rect 20138 5908 20174 5934
rect 20380 5908 20416 5934
rect 20474 5908 20510 5934
rect 20716 5908 20752 5934
rect 20810 5908 20846 5934
rect 21052 5908 21088 5934
rect 21146 5908 21182 5934
rect 21388 5908 21424 5934
rect 21482 5908 21518 5934
rect 21724 5908 21760 5934
rect 21818 5908 21854 5934
rect 29302 5908 29338 5934
rect 29396 5908 29432 5934
rect 29638 5908 29674 5934
rect 29732 5908 29768 5934
rect 29974 5908 30010 5934
rect 30068 5908 30104 5934
rect 30310 5908 30346 5934
rect 30404 5908 30440 5934
rect 30646 5908 30682 5934
rect 30740 5908 30776 5934
rect 30982 5908 31018 5934
rect 31076 5908 31112 5934
rect -4464 5862 -4428 5884
rect -4370 5862 -4334 5884
rect -4128 5862 -4092 5884
rect -4034 5862 -3998 5884
rect -3792 5862 -3756 5884
rect -3698 5862 -3662 5884
rect -3456 5862 -3420 5884
rect -3362 5862 -3326 5884
rect -3120 5862 -3084 5884
rect -3026 5862 -2990 5884
rect -2784 5862 -2748 5884
rect -2690 5862 -2654 5884
rect -4479 5846 -4319 5862
rect -4479 5812 -4463 5846
rect -4429 5812 -4369 5846
rect -4335 5812 -4319 5846
rect -4479 5796 -4319 5812
rect -4143 5846 -3983 5862
rect -4143 5812 -4127 5846
rect -4093 5812 -4033 5846
rect -3999 5812 -3983 5846
rect -4143 5796 -3983 5812
rect -3807 5846 -3647 5862
rect -3807 5812 -3791 5846
rect -3757 5812 -3697 5846
rect -3663 5812 -3647 5846
rect -3807 5796 -3647 5812
rect -3471 5846 -3311 5862
rect -3471 5812 -3455 5846
rect -3421 5812 -3361 5846
rect -3327 5812 -3311 5846
rect -3471 5796 -3311 5812
rect -3135 5846 -2975 5862
rect -3135 5812 -3119 5846
rect -3085 5812 -3025 5846
rect -2991 5812 -2975 5846
rect -3135 5796 -2975 5812
rect -2799 5846 -2639 5862
rect -2799 5812 -2783 5846
rect -2749 5812 -2689 5846
rect -2655 5812 -2639 5846
rect -2799 5796 -2639 5812
<< polycont >>
rect -4652 8407 -4614 8441
rect -4524 8407 -4486 8441
rect -4248 8407 -4210 8441
rect -4120 8407 -4082 8441
rect -3844 8407 -3806 8441
rect -3716 8407 -3678 8441
rect -3440 8407 -3402 8441
rect -3312 8407 -3274 8441
rect -3036 8407 -2998 8441
rect -2908 8407 -2870 8441
rect -2632 8407 -2594 8441
rect -2504 8407 -2466 8441
rect -4652 7279 -4614 7313
rect -4524 7279 -4486 7313
rect -4248 7279 -4210 7313
rect -4120 7279 -4082 7313
rect -3844 7279 -3806 7313
rect -3716 7279 -3678 7313
rect -3440 7279 -3402 7313
rect -3312 7279 -3274 7313
rect -3036 7279 -2998 7313
rect -2908 7279 -2870 7313
rect -2632 7279 -2594 7313
rect 746 7329 784 7363
rect 874 7329 912 7363
rect 1150 7329 1188 7363
rect 1278 7329 1316 7363
rect 1554 7329 1592 7363
rect 1682 7329 1720 7363
rect 1958 7329 1996 7363
rect 2086 7329 2124 7363
rect 2362 7329 2400 7363
rect 2490 7329 2528 7363
rect 2766 7329 2804 7363
rect 2894 7329 2932 7363
rect 7116 7329 7154 7363
rect 7244 7329 7282 7363
rect 7520 7329 7558 7363
rect 7648 7329 7686 7363
rect 7924 7329 7962 7363
rect 8052 7329 8090 7363
rect 8328 7329 8366 7363
rect 8456 7329 8494 7363
rect 8732 7329 8770 7363
rect 8860 7329 8898 7363
rect 9136 7329 9174 7363
rect 9264 7329 9302 7363
rect 13486 7329 13524 7363
rect 13614 7329 13652 7363
rect 13890 7329 13928 7363
rect 14018 7329 14056 7363
rect 14294 7329 14332 7363
rect 14422 7329 14460 7363
rect 14698 7329 14736 7363
rect 14826 7329 14864 7363
rect 15102 7329 15140 7363
rect 15230 7329 15268 7363
rect 15506 7329 15544 7363
rect 15634 7329 15672 7363
rect 19856 7329 19894 7363
rect 19984 7329 20022 7363
rect 20260 7329 20298 7363
rect 20388 7329 20426 7363
rect 20664 7329 20702 7363
rect 20792 7329 20830 7363
rect 21068 7329 21106 7363
rect 21196 7329 21234 7363
rect 21472 7329 21510 7363
rect 21600 7329 21638 7363
rect 21876 7329 21914 7363
rect 22004 7329 22042 7363
rect 29114 7329 29152 7363
rect 29242 7329 29280 7363
rect 29518 7329 29556 7363
rect 29646 7329 29684 7363
rect 29922 7329 29960 7363
rect 30050 7329 30088 7363
rect 30326 7329 30364 7363
rect 30454 7329 30492 7363
rect 30730 7329 30768 7363
rect 30858 7329 30896 7363
rect 31134 7329 31172 7363
rect 31262 7329 31300 7363
rect -2504 7279 -2466 7313
rect 935 6972 969 7006
rect 1029 6972 1063 7006
rect -4463 6922 -4429 6956
rect -4369 6922 -4335 6956
rect -4127 6922 -4093 6956
rect -4033 6922 -3999 6956
rect -3791 6922 -3757 6956
rect -3697 6922 -3663 6956
rect -3455 6922 -3421 6956
rect -3361 6922 -3327 6956
rect -3119 6922 -3085 6956
rect -3025 6922 -2991 6956
rect 1271 6972 1305 7006
rect 1365 6972 1399 7006
rect 1607 6972 1641 7006
rect 1701 6972 1735 7006
rect 1943 6972 1977 7006
rect 2037 6972 2071 7006
rect 2279 6972 2313 7006
rect 2373 6972 2407 7006
rect 2615 6972 2649 7006
rect 2709 6972 2743 7006
rect 7305 6972 7339 7006
rect 7399 6972 7433 7006
rect 7641 6972 7675 7006
rect 7735 6972 7769 7006
rect 7977 6972 8011 7006
rect 8071 6972 8105 7006
rect 8313 6972 8347 7006
rect 8407 6972 8441 7006
rect 8649 6972 8683 7006
rect 8743 6972 8777 7006
rect 8985 6972 9019 7006
rect 9079 6972 9113 7006
rect 13675 6972 13709 7006
rect 13769 6972 13803 7006
rect 14011 6972 14045 7006
rect 14105 6972 14139 7006
rect 14347 6972 14381 7006
rect 14441 6972 14475 7006
rect 14683 6972 14717 7006
rect 14777 6972 14811 7006
rect 15019 6972 15053 7006
rect 15113 6972 15147 7006
rect 15355 6972 15389 7006
rect 15449 6972 15483 7006
rect 20045 6972 20079 7006
rect 20139 6972 20173 7006
rect 20381 6972 20415 7006
rect 20475 6972 20509 7006
rect 20717 6972 20751 7006
rect 20811 6972 20845 7006
rect 21053 6972 21087 7006
rect 21147 6972 21181 7006
rect 21389 6972 21423 7006
rect 21483 6972 21517 7006
rect 21725 6972 21759 7006
rect 21819 6972 21853 7006
rect 29303 6972 29337 7006
rect 29397 6972 29431 7006
rect 29639 6972 29673 7006
rect 29733 6972 29767 7006
rect 29975 6972 30009 7006
rect 30069 6972 30103 7006
rect 30311 6972 30345 7006
rect 30405 6972 30439 7006
rect 30647 6972 30681 7006
rect 30741 6972 30775 7006
rect 30983 6972 31017 7006
rect 31077 6972 31111 7006
rect -2783 6922 -2749 6956
rect -2689 6922 -2655 6956
rect -4463 5812 -4429 5846
rect -4369 5812 -4335 5846
rect -4127 5812 -4093 5846
rect -4033 5812 -3999 5846
rect -3791 5812 -3757 5846
rect -3697 5812 -3663 5846
rect -3455 5812 -3421 5846
rect -3361 5812 -3327 5846
rect -3119 5812 -3085 5846
rect -3025 5812 -2991 5846
rect -2783 5812 -2749 5846
rect -2689 5812 -2655 5846
<< locali >>
rect -4668 8407 -4652 8441
rect -4614 8407 -4598 8441
rect -4540 8407 -4524 8441
rect -4486 8407 -4470 8441
rect -4264 8407 -4248 8441
rect -4210 8407 -4194 8441
rect -4136 8407 -4120 8441
rect -4082 8407 -4066 8441
rect -3860 8407 -3844 8441
rect -3806 8407 -3790 8441
rect -3732 8407 -3716 8441
rect -3678 8407 -3662 8441
rect -3456 8407 -3440 8441
rect -3402 8407 -3386 8441
rect -3328 8407 -3312 8441
rect -3274 8407 -3258 8441
rect -3052 8407 -3036 8441
rect -2998 8407 -2982 8441
rect -2924 8407 -2908 8441
rect -2870 8407 -2854 8441
rect -2648 8407 -2632 8441
rect -2594 8407 -2578 8441
rect -2520 8407 -2504 8441
rect -2466 8407 -2450 8441
rect 610 8398 644 8414
rect -4788 8348 -4754 8364
rect -4788 7356 -4754 7372
rect -4714 8348 -4680 8364
rect -4714 7356 -4680 7372
rect -4586 8348 -4552 8364
rect -4586 7356 -4552 7372
rect -4458 8348 -4424 8364
rect -4458 7356 -4424 7372
rect -4384 8348 -4350 8364
rect -4384 7356 -4350 7372
rect -4310 8348 -4276 8364
rect -4310 7356 -4276 7372
rect -4182 8348 -4148 8364
rect -4182 7356 -4148 7372
rect -4054 8348 -4020 8364
rect -4054 7356 -4020 7372
rect -3980 8348 -3946 8364
rect -3980 7356 -3946 7372
rect -3906 8348 -3872 8364
rect -3906 7356 -3872 7372
rect -3778 8348 -3744 8364
rect -3778 7356 -3744 7372
rect -3650 8348 -3616 8364
rect -3650 7356 -3616 7372
rect -3576 8348 -3542 8364
rect -3576 7356 -3542 7372
rect -3502 8348 -3468 8364
rect -3502 7356 -3468 7372
rect -3374 8348 -3340 8364
rect -3374 7356 -3340 7372
rect -3246 8348 -3212 8364
rect -3246 7356 -3212 7372
rect -3172 8348 -3138 8364
rect -3172 7356 -3138 7372
rect -3098 8348 -3064 8364
rect -3098 7356 -3064 7372
rect -2970 8348 -2936 8364
rect -2970 7356 -2936 7372
rect -2842 8348 -2808 8364
rect -2842 7356 -2808 7372
rect -2768 8348 -2734 8364
rect -2768 7356 -2734 7372
rect -2694 8348 -2660 8364
rect -2694 7356 -2660 7372
rect -2566 8348 -2532 8364
rect -2566 7356 -2532 7372
rect -2438 8348 -2404 8364
rect -2438 7356 -2404 7372
rect -2364 8348 -2330 8364
rect 610 7406 644 7422
rect 684 8398 718 8414
rect 684 7406 718 7422
rect 812 8398 846 8414
rect 812 7406 846 7422
rect 940 8398 974 8414
rect 940 7406 974 7422
rect 1014 8398 1048 8414
rect 1014 7406 1048 7422
rect 1088 8398 1122 8414
rect 1088 7406 1122 7422
rect 1216 8398 1250 8414
rect 1216 7406 1250 7422
rect 1344 8398 1378 8414
rect 1344 7406 1378 7422
rect 1418 8398 1452 8414
rect 1418 7406 1452 7422
rect 1492 8398 1526 8414
rect 1492 7406 1526 7422
rect 1620 8398 1654 8414
rect 1620 7406 1654 7422
rect 1748 8398 1782 8414
rect 1748 7406 1782 7422
rect 1822 8398 1856 8414
rect 1822 7406 1856 7422
rect 1896 8398 1930 8414
rect 1896 7406 1930 7422
rect 2024 8398 2058 8414
rect 2024 7406 2058 7422
rect 2152 8398 2186 8414
rect 2152 7406 2186 7422
rect 2226 8398 2260 8414
rect 2226 7406 2260 7422
rect 2300 8398 2334 8414
rect 2300 7406 2334 7422
rect 2428 8398 2462 8414
rect 2428 7406 2462 7422
rect 2556 8398 2590 8414
rect 2556 7406 2590 7422
rect 2630 8398 2664 8414
rect 2630 7406 2664 7422
rect 2704 8398 2738 8414
rect 2704 7406 2738 7422
rect 2832 8398 2866 8414
rect 2832 7406 2866 7422
rect 2960 8398 2994 8414
rect 2960 7406 2994 7422
rect 3034 8398 3068 8414
rect 3034 7406 3068 7422
rect 6980 8398 7014 8414
rect 6980 7406 7014 7422
rect 7054 8398 7088 8414
rect 7054 7406 7088 7422
rect 7182 8398 7216 8414
rect 7182 7406 7216 7422
rect 7310 8398 7344 8414
rect 7310 7406 7344 7422
rect 7384 8398 7418 8414
rect 7384 7406 7418 7422
rect 7458 8398 7492 8414
rect 7458 7406 7492 7422
rect 7586 8398 7620 8414
rect 7586 7406 7620 7422
rect 7714 8398 7748 8414
rect 7714 7406 7748 7422
rect 7788 8398 7822 8414
rect 7788 7406 7822 7422
rect 7862 8398 7896 8414
rect 7862 7406 7896 7422
rect 7990 8398 8024 8414
rect 7990 7406 8024 7422
rect 8118 8398 8152 8414
rect 8118 7406 8152 7422
rect 8192 8398 8226 8414
rect 8192 7406 8226 7422
rect 8266 8398 8300 8414
rect 8266 7406 8300 7422
rect 8394 8398 8428 8414
rect 8394 7406 8428 7422
rect 8522 8398 8556 8414
rect 8522 7406 8556 7422
rect 8596 8398 8630 8414
rect 8596 7406 8630 7422
rect 8670 8398 8704 8414
rect 8670 7406 8704 7422
rect 8798 8398 8832 8414
rect 8798 7406 8832 7422
rect 8926 8398 8960 8414
rect 8926 7406 8960 7422
rect 9000 8398 9034 8414
rect 9000 7406 9034 7422
rect 9074 8398 9108 8414
rect 9074 7406 9108 7422
rect 9202 8398 9236 8414
rect 9202 7406 9236 7422
rect 9330 8398 9364 8414
rect 9330 7406 9364 7422
rect 9404 8398 9438 8414
rect 9404 7406 9438 7422
rect 13350 8398 13384 8414
rect 13350 7406 13384 7422
rect 13424 8398 13458 8414
rect 13424 7406 13458 7422
rect 13552 8398 13586 8414
rect 13552 7406 13586 7422
rect 13680 8398 13714 8414
rect 13680 7406 13714 7422
rect 13754 8398 13788 8414
rect 13754 7406 13788 7422
rect 13828 8398 13862 8414
rect 13828 7406 13862 7422
rect 13956 8398 13990 8414
rect 13956 7406 13990 7422
rect 14084 8398 14118 8414
rect 14084 7406 14118 7422
rect 14158 8398 14192 8414
rect 14158 7406 14192 7422
rect 14232 8398 14266 8414
rect 14232 7406 14266 7422
rect 14360 8398 14394 8414
rect 14360 7406 14394 7422
rect 14488 8398 14522 8414
rect 14488 7406 14522 7422
rect 14562 8398 14596 8414
rect 14562 7406 14596 7422
rect 14636 8398 14670 8414
rect 14636 7406 14670 7422
rect 14764 8398 14798 8414
rect 14764 7406 14798 7422
rect 14892 8398 14926 8414
rect 14892 7406 14926 7422
rect 14966 8398 15000 8414
rect 14966 7406 15000 7422
rect 15040 8398 15074 8414
rect 15040 7406 15074 7422
rect 15168 8398 15202 8414
rect 15168 7406 15202 7422
rect 15296 8398 15330 8414
rect 15296 7406 15330 7422
rect 15370 8398 15404 8414
rect 15370 7406 15404 7422
rect 15444 8398 15478 8414
rect 15444 7406 15478 7422
rect 15572 8398 15606 8414
rect 15572 7406 15606 7422
rect 15700 8398 15734 8414
rect 15700 7406 15734 7422
rect 15774 8398 15808 8414
rect 15774 7406 15808 7422
rect 19720 8398 19754 8414
rect 19720 7406 19754 7422
rect 19794 8398 19828 8414
rect 19794 7406 19828 7422
rect 19922 8398 19956 8414
rect 19922 7406 19956 7422
rect 20050 8398 20084 8414
rect 20050 7406 20084 7422
rect 20124 8398 20158 8414
rect 20124 7406 20158 7422
rect 20198 8398 20232 8414
rect 20198 7406 20232 7422
rect 20326 8398 20360 8414
rect 20326 7406 20360 7422
rect 20454 8398 20488 8414
rect 20454 7406 20488 7422
rect 20528 8398 20562 8414
rect 20528 7406 20562 7422
rect 20602 8398 20636 8414
rect 20602 7406 20636 7422
rect 20730 8398 20764 8414
rect 20730 7406 20764 7422
rect 20858 8398 20892 8414
rect 20858 7406 20892 7422
rect 20932 8398 20966 8414
rect 20932 7406 20966 7422
rect 21006 8398 21040 8414
rect 21006 7406 21040 7422
rect 21134 8398 21168 8414
rect 21134 7406 21168 7422
rect 21262 8398 21296 8414
rect 21262 7406 21296 7422
rect 21336 8398 21370 8414
rect 21336 7406 21370 7422
rect 21410 8398 21444 8414
rect 21410 7406 21444 7422
rect 21538 8398 21572 8414
rect 21538 7406 21572 7422
rect 21666 8398 21700 8414
rect 21666 7406 21700 7422
rect 21740 8398 21774 8414
rect 21740 7406 21774 7422
rect 21814 8398 21848 8414
rect 21814 7406 21848 7422
rect 21942 8398 21976 8414
rect 21942 7406 21976 7422
rect 22070 8398 22104 8414
rect 22070 7406 22104 7422
rect 22144 8398 22178 8414
rect 22144 7406 22178 7422
rect 28978 8398 29012 8414
rect 28978 7406 29012 7422
rect 29052 8398 29086 8414
rect 29052 7406 29086 7422
rect 29180 8398 29214 8414
rect 29180 7406 29214 7422
rect 29308 8398 29342 8414
rect 29308 7406 29342 7422
rect 29382 8398 29416 8414
rect 29382 7406 29416 7422
rect 29456 8398 29490 8414
rect 29456 7406 29490 7422
rect 29584 8398 29618 8414
rect 29584 7406 29618 7422
rect 29712 8398 29746 8414
rect 29712 7406 29746 7422
rect 29786 8398 29820 8414
rect 29786 7406 29820 7422
rect 29860 8398 29894 8414
rect 29860 7406 29894 7422
rect 29988 8398 30022 8414
rect 29988 7406 30022 7422
rect 30116 8398 30150 8414
rect 30116 7406 30150 7422
rect 30190 8398 30224 8414
rect 30190 7406 30224 7422
rect 30264 8398 30298 8414
rect 30264 7406 30298 7422
rect 30392 8398 30426 8414
rect 30392 7406 30426 7422
rect 30520 8398 30554 8414
rect 30520 7406 30554 7422
rect 30594 8398 30628 8414
rect 30594 7406 30628 7422
rect 30668 8398 30702 8414
rect 30668 7406 30702 7422
rect 30796 8398 30830 8414
rect 30796 7406 30830 7422
rect 30924 8398 30958 8414
rect 30924 7406 30958 7422
rect 30998 8398 31032 8414
rect 30998 7406 31032 7422
rect 31072 8398 31106 8414
rect 31072 7406 31106 7422
rect 31200 8398 31234 8414
rect 31200 7406 31234 7422
rect 31328 8398 31362 8414
rect 31328 7406 31362 7422
rect 31402 8398 31436 8414
rect 31402 7406 31436 7422
rect -2364 7356 -2330 7372
rect 730 7329 746 7363
rect 784 7329 800 7363
rect 858 7329 874 7363
rect 912 7329 928 7363
rect 1134 7329 1150 7363
rect 1188 7329 1204 7363
rect 1262 7329 1278 7363
rect 1316 7329 1332 7363
rect 1538 7329 1554 7363
rect 1592 7329 1608 7363
rect 1666 7329 1682 7363
rect 1720 7329 1736 7363
rect 1942 7329 1958 7363
rect 1996 7329 2012 7363
rect 2070 7329 2086 7363
rect 2124 7329 2140 7363
rect 2346 7329 2362 7363
rect 2400 7329 2416 7363
rect 2474 7329 2490 7363
rect 2528 7329 2544 7363
rect 2750 7329 2766 7363
rect 2804 7329 2820 7363
rect 2878 7329 2894 7363
rect 2932 7329 2948 7363
rect 7100 7329 7116 7363
rect 7154 7329 7170 7363
rect 7228 7329 7244 7363
rect 7282 7329 7298 7363
rect 7504 7329 7520 7363
rect 7558 7329 7574 7363
rect 7632 7329 7648 7363
rect 7686 7329 7702 7363
rect 7908 7329 7924 7363
rect 7962 7329 7978 7363
rect 8036 7329 8052 7363
rect 8090 7329 8106 7363
rect 8312 7329 8328 7363
rect 8366 7329 8382 7363
rect 8440 7329 8456 7363
rect 8494 7329 8510 7363
rect 8716 7329 8732 7363
rect 8770 7329 8786 7363
rect 8844 7329 8860 7363
rect 8898 7329 8914 7363
rect 9120 7329 9136 7363
rect 9174 7329 9190 7363
rect 9248 7329 9264 7363
rect 9302 7329 9318 7363
rect 13470 7329 13486 7363
rect 13524 7329 13540 7363
rect 13598 7329 13614 7363
rect 13652 7329 13668 7363
rect 13874 7329 13890 7363
rect 13928 7329 13944 7363
rect 14002 7329 14018 7363
rect 14056 7329 14072 7363
rect 14278 7329 14294 7363
rect 14332 7329 14348 7363
rect 14406 7329 14422 7363
rect 14460 7329 14476 7363
rect 14682 7329 14698 7363
rect 14736 7329 14752 7363
rect 14810 7329 14826 7363
rect 14864 7329 14880 7363
rect 15086 7329 15102 7363
rect 15140 7329 15156 7363
rect 15214 7329 15230 7363
rect 15268 7329 15284 7363
rect 15490 7329 15506 7363
rect 15544 7329 15560 7363
rect 15618 7329 15634 7363
rect 15672 7329 15688 7363
rect 19840 7329 19856 7363
rect 19894 7329 19910 7363
rect 19968 7329 19984 7363
rect 20022 7329 20038 7363
rect 20244 7329 20260 7363
rect 20298 7329 20314 7363
rect 20372 7329 20388 7363
rect 20426 7329 20442 7363
rect 20648 7329 20664 7363
rect 20702 7329 20718 7363
rect 20776 7329 20792 7363
rect 20830 7329 20846 7363
rect 21052 7329 21068 7363
rect 21106 7329 21122 7363
rect 21180 7329 21196 7363
rect 21234 7329 21250 7363
rect 21456 7329 21472 7363
rect 21510 7329 21526 7363
rect 21584 7329 21600 7363
rect 21638 7329 21654 7363
rect 21860 7329 21876 7363
rect 21914 7329 21930 7363
rect 21988 7329 22004 7363
rect 22042 7329 22058 7363
rect 29098 7329 29114 7363
rect 29152 7329 29168 7363
rect 29226 7329 29242 7363
rect 29280 7329 29296 7363
rect 29502 7329 29518 7363
rect 29556 7329 29572 7363
rect 29630 7329 29646 7363
rect 29684 7329 29700 7363
rect 29906 7329 29922 7363
rect 29960 7329 29976 7363
rect 30034 7329 30050 7363
rect 30088 7329 30104 7363
rect 30310 7329 30326 7363
rect 30364 7329 30380 7363
rect 30438 7329 30454 7363
rect 30492 7329 30508 7363
rect 30714 7329 30730 7363
rect 30768 7329 30784 7363
rect 30842 7329 30858 7363
rect 30896 7329 30912 7363
rect 31118 7329 31134 7363
rect 31172 7329 31188 7363
rect 31246 7329 31262 7363
rect 31300 7329 31316 7363
rect -4668 7279 -4652 7313
rect -4614 7279 -4598 7313
rect -4540 7279 -4524 7313
rect -4486 7279 -4470 7313
rect -4264 7279 -4248 7313
rect -4210 7279 -4194 7313
rect -4136 7279 -4120 7313
rect -4082 7279 -4066 7313
rect -3860 7279 -3844 7313
rect -3806 7279 -3790 7313
rect -3732 7279 -3716 7313
rect -3678 7279 -3662 7313
rect -3456 7279 -3440 7313
rect -3402 7279 -3386 7313
rect -3328 7279 -3312 7313
rect -3274 7279 -3258 7313
rect -3052 7279 -3036 7313
rect -2998 7279 -2982 7313
rect -2924 7279 -2908 7313
rect -2870 7279 -2854 7313
rect -2648 7279 -2632 7313
rect -2594 7279 -2578 7313
rect -2520 7279 -2504 7313
rect -2466 7279 -2450 7313
rect 919 6972 935 7006
rect 969 6972 1029 7006
rect 1063 6972 1079 7006
rect 1255 6972 1271 7006
rect 1305 6972 1365 7006
rect 1399 6972 1415 7006
rect 1591 6972 1607 7006
rect 1641 6972 1701 7006
rect 1735 6972 1751 7006
rect 1927 6972 1943 7006
rect 1977 6972 2037 7006
rect 2071 6972 2087 7006
rect 2263 6972 2279 7006
rect 2313 6972 2373 7006
rect 2407 6972 2423 7006
rect 2599 6972 2615 7006
rect 2649 6972 2709 7006
rect 2743 6972 2759 7006
rect 7289 6972 7305 7006
rect 7339 6972 7399 7006
rect 7433 6972 7449 7006
rect 7625 6972 7641 7006
rect 7675 6972 7735 7006
rect 7769 6972 7785 7006
rect 7961 6972 7977 7006
rect 8011 6972 8071 7006
rect 8105 6972 8121 7006
rect 8297 6972 8313 7006
rect 8347 6972 8407 7006
rect 8441 6972 8457 7006
rect 8633 6972 8649 7006
rect 8683 6972 8743 7006
rect 8777 6972 8793 7006
rect 8969 6972 8985 7006
rect 9019 6972 9079 7006
rect 9113 6972 9129 7006
rect 13659 6972 13675 7006
rect 13709 6972 13769 7006
rect 13803 6972 13819 7006
rect 13995 6972 14011 7006
rect 14045 6972 14105 7006
rect 14139 6972 14155 7006
rect 14331 6972 14347 7006
rect 14381 6972 14441 7006
rect 14475 6972 14491 7006
rect 14667 6972 14683 7006
rect 14717 6972 14777 7006
rect 14811 6972 14827 7006
rect 15003 6972 15019 7006
rect 15053 6972 15113 7006
rect 15147 6972 15163 7006
rect 15339 6972 15355 7006
rect 15389 6972 15449 7006
rect 15483 6972 15499 7006
rect 20029 6972 20045 7006
rect 20079 6972 20139 7006
rect 20173 6972 20189 7006
rect 20365 6972 20381 7006
rect 20415 6972 20475 7006
rect 20509 6972 20525 7006
rect 20701 6972 20717 7006
rect 20751 6972 20811 7006
rect 20845 6972 20861 7006
rect 21037 6972 21053 7006
rect 21087 6972 21147 7006
rect 21181 6972 21197 7006
rect 21373 6972 21389 7006
rect 21423 6972 21483 7006
rect 21517 6972 21533 7006
rect 21709 6972 21725 7006
rect 21759 6972 21819 7006
rect 21853 6972 21869 7006
rect 29287 6972 29303 7006
rect 29337 6972 29397 7006
rect 29431 6972 29447 7006
rect 29623 6972 29639 7006
rect 29673 6972 29733 7006
rect 29767 6972 29783 7006
rect 29959 6972 29975 7006
rect 30009 6972 30069 7006
rect 30103 6972 30119 7006
rect 30295 6972 30311 7006
rect 30345 6972 30405 7006
rect 30439 6972 30455 7006
rect 30631 6972 30647 7006
rect 30681 6972 30741 7006
rect 30775 6972 30791 7006
rect 30967 6972 30983 7006
rect 31017 6972 31077 7006
rect 31111 6972 31127 7006
rect -4479 6922 -4463 6956
rect -4429 6922 -4369 6956
rect -4335 6922 -4319 6956
rect -4143 6922 -4127 6956
rect -4093 6922 -4033 6956
rect -3999 6922 -3983 6956
rect -3807 6922 -3791 6956
rect -3757 6922 -3697 6956
rect -3663 6922 -3647 6956
rect -3471 6922 -3455 6956
rect -3421 6922 -3361 6956
rect -3327 6922 -3311 6956
rect -3135 6922 -3119 6956
rect -3085 6922 -3025 6956
rect -2991 6922 -2975 6956
rect -2799 6922 -2783 6956
rect -2749 6922 -2689 6956
rect -2655 6922 -2639 6956
rect -4584 6872 -4550 6888
rect -4584 5880 -4550 5896
rect -4510 6872 -4476 6888
rect -4510 5880 -4476 5896
rect -4416 6872 -4382 6888
rect -4416 5880 -4382 5896
rect -4322 6872 -4288 6888
rect -4322 5880 -4288 5896
rect -4248 6872 -4214 6888
rect -4248 5880 -4214 5896
rect -4174 6872 -4140 6888
rect -4174 5880 -4140 5896
rect -4080 6872 -4046 6888
rect -4080 5880 -4046 5896
rect -3986 6872 -3952 6888
rect -3986 5880 -3952 5896
rect -3912 6872 -3878 6888
rect -3912 5880 -3878 5896
rect -3838 6872 -3804 6888
rect -3838 5880 -3804 5896
rect -3744 6872 -3710 6888
rect -3744 5880 -3710 5896
rect -3650 6872 -3616 6888
rect -3650 5880 -3616 5896
rect -3576 6872 -3542 6888
rect -3576 5880 -3542 5896
rect -3502 6872 -3468 6888
rect -3502 5880 -3468 5896
rect -3408 6872 -3374 6888
rect -3408 5880 -3374 5896
rect -3314 6872 -3280 6888
rect -3314 5880 -3280 5896
rect -3240 6872 -3206 6888
rect -3240 5880 -3206 5896
rect -3166 6872 -3132 6888
rect -3166 5880 -3132 5896
rect -3072 6872 -3038 6888
rect -3072 5880 -3038 5896
rect -2978 6872 -2944 6888
rect -2978 5880 -2944 5896
rect -2904 6872 -2870 6888
rect -2904 5880 -2870 5896
rect -2830 6872 -2796 6888
rect -2830 5880 -2796 5896
rect -2736 6872 -2702 6888
rect -2736 5880 -2702 5896
rect -2642 6872 -2608 6888
rect -2642 5880 -2608 5896
rect -2568 6872 -2534 6888
rect 814 6880 848 6938
rect 814 6812 848 6846
rect 814 6744 848 6778
rect 814 6676 848 6710
rect 814 6634 848 6642
rect 814 5930 848 5946
rect 888 6922 922 6938
rect 888 5930 922 5946
rect 982 6922 1016 6938
rect 982 5930 1016 5946
rect 1076 6922 1110 6938
rect 1076 5930 1110 5946
rect 1150 6906 1184 6938
rect 1150 6838 1184 6872
rect 1150 6770 1184 6804
rect 1150 6702 1184 6736
rect 1150 6634 1184 6668
rect 1150 5930 1184 5946
rect 1224 6922 1258 6938
rect 1224 5930 1258 5946
rect 1318 6922 1352 6938
rect 1318 5930 1352 5946
rect 1412 6922 1446 6938
rect 1412 5930 1446 5946
rect 1486 6906 1520 6938
rect 1486 6838 1520 6872
rect 1486 6770 1520 6804
rect 1486 6702 1520 6736
rect 1486 6634 1520 6668
rect 1486 5930 1520 5946
rect 1560 6922 1594 6938
rect 1560 5930 1594 5946
rect 1654 6922 1688 6938
rect 1654 5930 1688 5946
rect 1748 6922 1782 6938
rect 1748 5930 1782 5946
rect 1822 6906 1856 6938
rect 1822 6838 1856 6872
rect 1822 6770 1856 6804
rect 1822 6702 1856 6736
rect 1822 6634 1856 6668
rect 1822 5930 1856 5946
rect 1896 6922 1930 6938
rect 1896 5930 1930 5946
rect 1990 6922 2024 6938
rect 1990 5930 2024 5946
rect 2084 6922 2118 6938
rect 2084 5930 2118 5946
rect 2158 6906 2192 6938
rect 2158 6838 2192 6872
rect 2158 6770 2192 6804
rect 2158 6702 2192 6736
rect 2158 6634 2192 6668
rect 2158 5930 2192 5946
rect 2232 6922 2266 6938
rect 2232 5930 2266 5946
rect 2326 6922 2360 6938
rect 2326 5930 2360 5946
rect 2420 6922 2454 6938
rect 2420 5930 2454 5946
rect 2494 6906 2528 6938
rect 2494 6838 2528 6872
rect 2494 6770 2528 6804
rect 2494 6702 2528 6736
rect 2494 6634 2528 6668
rect 2494 5930 2528 5946
rect 2568 6922 2602 6938
rect 2568 5930 2602 5946
rect 2662 6922 2696 6938
rect 2662 5930 2696 5946
rect 2756 6922 2790 6938
rect 2756 5930 2790 5946
rect 2830 6906 2864 6938
rect 2830 6838 2864 6872
rect 2830 6770 2864 6804
rect 2830 6702 2864 6736
rect 2830 6634 2864 6668
rect 2830 5930 2864 5946
rect 7184 6880 7218 6938
rect 7184 6812 7218 6846
rect 7184 6744 7218 6778
rect 7184 6676 7218 6710
rect 7184 6634 7218 6642
rect 7184 5930 7218 5946
rect 7258 6922 7292 6938
rect 7258 5930 7292 5946
rect 7352 6922 7386 6938
rect 7352 5930 7386 5946
rect 7446 6922 7480 6938
rect 7446 5930 7480 5946
rect 7520 6906 7554 6938
rect 7520 6838 7554 6872
rect 7520 6770 7554 6804
rect 7520 6702 7554 6736
rect 7520 6634 7554 6668
rect 7520 5930 7554 5946
rect 7594 6922 7628 6938
rect 7594 5930 7628 5946
rect 7688 6922 7722 6938
rect 7688 5930 7722 5946
rect 7782 6922 7816 6938
rect 7782 5930 7816 5946
rect 7856 6906 7890 6938
rect 7856 6838 7890 6872
rect 7856 6770 7890 6804
rect 7856 6702 7890 6736
rect 7856 6634 7890 6668
rect 7856 5930 7890 5946
rect 7930 6922 7964 6938
rect 7930 5930 7964 5946
rect 8024 6922 8058 6938
rect 8024 5930 8058 5946
rect 8118 6922 8152 6938
rect 8118 5930 8152 5946
rect 8192 6906 8226 6938
rect 8192 6838 8226 6872
rect 8192 6770 8226 6804
rect 8192 6702 8226 6736
rect 8192 6634 8226 6668
rect 8192 5930 8226 5946
rect 8266 6922 8300 6938
rect 8266 5930 8300 5946
rect 8360 6922 8394 6938
rect 8360 5930 8394 5946
rect 8454 6922 8488 6938
rect 8454 5930 8488 5946
rect 8528 6906 8562 6938
rect 8528 6838 8562 6872
rect 8528 6770 8562 6804
rect 8528 6702 8562 6736
rect 8528 6634 8562 6668
rect 8528 5930 8562 5946
rect 8602 6922 8636 6938
rect 8602 5930 8636 5946
rect 8696 6922 8730 6938
rect 8696 5930 8730 5946
rect 8790 6922 8824 6938
rect 8790 5930 8824 5946
rect 8864 6906 8898 6938
rect 8864 6838 8898 6872
rect 8864 6770 8898 6804
rect 8864 6702 8898 6736
rect 8864 6634 8898 6668
rect 8864 5930 8898 5946
rect 8938 6922 8972 6938
rect 8938 5930 8972 5946
rect 9032 6922 9066 6938
rect 9032 5930 9066 5946
rect 9126 6922 9160 6938
rect 9126 5930 9160 5946
rect 9200 6906 9234 6938
rect 9200 6838 9234 6872
rect 9200 6770 9234 6804
rect 9200 6702 9234 6736
rect 9200 6634 9234 6668
rect 9200 5930 9234 5946
rect 13554 6880 13588 6938
rect 13554 6812 13588 6846
rect 13554 6744 13588 6778
rect 13554 6676 13588 6710
rect 13554 6634 13588 6642
rect 13554 5930 13588 5946
rect 13628 6922 13662 6938
rect 13628 5930 13662 5946
rect 13722 6922 13756 6938
rect 13722 5930 13756 5946
rect 13816 6922 13850 6938
rect 13816 5930 13850 5946
rect 13890 6906 13924 6938
rect 13890 6838 13924 6872
rect 13890 6770 13924 6804
rect 13890 6702 13924 6736
rect 13890 6634 13924 6668
rect 13890 5930 13924 5946
rect 13964 6922 13998 6938
rect 13964 5930 13998 5946
rect 14058 6922 14092 6938
rect 14058 5930 14092 5946
rect 14152 6922 14186 6938
rect 14152 5930 14186 5946
rect 14226 6906 14260 6938
rect 14226 6838 14260 6872
rect 14226 6770 14260 6804
rect 14226 6702 14260 6736
rect 14226 6634 14260 6668
rect 14226 5930 14260 5946
rect 14300 6922 14334 6938
rect 14300 5930 14334 5946
rect 14394 6922 14428 6938
rect 14394 5930 14428 5946
rect 14488 6922 14522 6938
rect 14488 5930 14522 5946
rect 14562 6906 14596 6938
rect 14562 6838 14596 6872
rect 14562 6770 14596 6804
rect 14562 6702 14596 6736
rect 14562 6634 14596 6668
rect 14562 5930 14596 5946
rect 14636 6922 14670 6938
rect 14636 5930 14670 5946
rect 14730 6922 14764 6938
rect 14730 5930 14764 5946
rect 14824 6922 14858 6938
rect 14824 5930 14858 5946
rect 14898 6906 14932 6938
rect 14898 6838 14932 6872
rect 14898 6770 14932 6804
rect 14898 6702 14932 6736
rect 14898 6634 14932 6668
rect 14898 5930 14932 5946
rect 14972 6922 15006 6938
rect 14972 5930 15006 5946
rect 15066 6922 15100 6938
rect 15066 5930 15100 5946
rect 15160 6922 15194 6938
rect 15160 5930 15194 5946
rect 15234 6906 15268 6938
rect 15234 6838 15268 6872
rect 15234 6770 15268 6804
rect 15234 6702 15268 6736
rect 15234 6634 15268 6668
rect 15234 5930 15268 5946
rect 15308 6922 15342 6938
rect 15308 5930 15342 5946
rect 15402 6922 15436 6938
rect 15402 5930 15436 5946
rect 15496 6922 15530 6938
rect 15496 5930 15530 5946
rect 15570 6906 15604 6938
rect 15570 6838 15604 6872
rect 15570 6770 15604 6804
rect 15570 6702 15604 6736
rect 15570 6634 15604 6668
rect 15570 5930 15604 5946
rect 19924 6880 19958 6938
rect 19924 6812 19958 6846
rect 19924 6744 19958 6778
rect 19924 6676 19958 6710
rect 19924 6634 19958 6642
rect 19924 5930 19958 5946
rect 19998 6922 20032 6938
rect 19998 5930 20032 5946
rect 20092 6922 20126 6938
rect 20092 5930 20126 5946
rect 20186 6922 20220 6938
rect 20186 5930 20220 5946
rect 20260 6906 20294 6938
rect 20260 6838 20294 6872
rect 20260 6770 20294 6804
rect 20260 6702 20294 6736
rect 20260 6634 20294 6668
rect 20260 5930 20294 5946
rect 20334 6922 20368 6938
rect 20334 5930 20368 5946
rect 20428 6922 20462 6938
rect 20428 5930 20462 5946
rect 20522 6922 20556 6938
rect 20522 5930 20556 5946
rect 20596 6906 20630 6938
rect 20596 6838 20630 6872
rect 20596 6770 20630 6804
rect 20596 6702 20630 6736
rect 20596 6634 20630 6668
rect 20596 5930 20630 5946
rect 20670 6922 20704 6938
rect 20670 5930 20704 5946
rect 20764 6922 20798 6938
rect 20764 5930 20798 5946
rect 20858 6922 20892 6938
rect 20858 5930 20892 5946
rect 20932 6906 20966 6938
rect 20932 6838 20966 6872
rect 20932 6770 20966 6804
rect 20932 6702 20966 6736
rect 20932 6634 20966 6668
rect 20932 5930 20966 5946
rect 21006 6922 21040 6938
rect 21006 5930 21040 5946
rect 21100 6922 21134 6938
rect 21100 5930 21134 5946
rect 21194 6922 21228 6938
rect 21194 5930 21228 5946
rect 21268 6906 21302 6938
rect 21268 6838 21302 6872
rect 21268 6770 21302 6804
rect 21268 6702 21302 6736
rect 21268 6634 21302 6668
rect 21268 5930 21302 5946
rect 21342 6922 21376 6938
rect 21342 5930 21376 5946
rect 21436 6922 21470 6938
rect 21436 5930 21470 5946
rect 21530 6922 21564 6938
rect 21530 5930 21564 5946
rect 21604 6906 21638 6938
rect 21604 6838 21638 6872
rect 21604 6770 21638 6804
rect 21604 6702 21638 6736
rect 21604 6634 21638 6668
rect 21604 5930 21638 5946
rect 21678 6922 21712 6938
rect 21678 5930 21712 5946
rect 21772 6922 21806 6938
rect 21772 5930 21806 5946
rect 21866 6922 21900 6938
rect 21866 5930 21900 5946
rect 21940 6906 21974 6938
rect 21940 6838 21974 6872
rect 21940 6770 21974 6804
rect 21940 6702 21974 6736
rect 21940 6634 21974 6668
rect 21940 5930 21974 5946
rect 29182 6880 29216 6938
rect 29182 6812 29216 6846
rect 29182 6744 29216 6778
rect 29182 6676 29216 6710
rect 29182 6634 29216 6642
rect 29182 5930 29216 5946
rect 29256 6922 29290 6938
rect 29256 5930 29290 5946
rect 29350 6922 29384 6938
rect 29350 5930 29384 5946
rect 29444 6922 29478 6938
rect 29444 5930 29478 5946
rect 29518 6906 29552 6938
rect 29518 6838 29552 6872
rect 29518 6770 29552 6804
rect 29518 6702 29552 6736
rect 29518 6634 29552 6668
rect 29518 5930 29552 5946
rect 29592 6922 29626 6938
rect 29592 5930 29626 5946
rect 29686 6922 29720 6938
rect 29686 5930 29720 5946
rect 29780 6922 29814 6938
rect 29780 5930 29814 5946
rect 29854 6906 29888 6938
rect 29854 6838 29888 6872
rect 29854 6770 29888 6804
rect 29854 6702 29888 6736
rect 29854 6634 29888 6668
rect 29854 5930 29888 5946
rect 29928 6922 29962 6938
rect 29928 5930 29962 5946
rect 30022 6922 30056 6938
rect 30022 5930 30056 5946
rect 30116 6922 30150 6938
rect 30116 5930 30150 5946
rect 30190 6906 30224 6938
rect 30190 6838 30224 6872
rect 30190 6770 30224 6804
rect 30190 6702 30224 6736
rect 30190 6634 30224 6668
rect 30190 5930 30224 5946
rect 30264 6922 30298 6938
rect 30264 5930 30298 5946
rect 30358 6922 30392 6938
rect 30358 5930 30392 5946
rect 30452 6922 30486 6938
rect 30452 5930 30486 5946
rect 30526 6906 30560 6938
rect 30526 6838 30560 6872
rect 30526 6770 30560 6804
rect 30526 6702 30560 6736
rect 30526 6634 30560 6668
rect 30526 5930 30560 5946
rect 30600 6922 30634 6938
rect 30600 5930 30634 5946
rect 30694 6922 30728 6938
rect 30694 5930 30728 5946
rect 30788 6922 30822 6938
rect 30788 5930 30822 5946
rect 30862 6906 30896 6938
rect 30862 6838 30896 6872
rect 30862 6770 30896 6804
rect 30862 6702 30896 6736
rect 30862 6634 30896 6668
rect 30862 5930 30896 5946
rect 30936 6922 30970 6938
rect 30936 5930 30970 5946
rect 31030 6922 31064 6938
rect 31030 5930 31064 5946
rect 31124 6922 31158 6938
rect 31124 5930 31158 5946
rect 31198 6906 31232 6938
rect 31198 6838 31232 6872
rect 31198 6770 31232 6804
rect 31198 6702 31232 6736
rect 31198 6634 31232 6668
rect 31198 5930 31232 5946
rect -2568 5880 -2534 5896
rect -4479 5812 -4463 5846
rect -4429 5812 -4369 5846
rect -4335 5812 -4319 5846
rect -4143 5812 -4127 5846
rect -4093 5812 -4033 5846
rect -3999 5812 -3983 5846
rect -3807 5812 -3791 5846
rect -3757 5812 -3697 5846
rect -3663 5812 -3647 5846
rect -3471 5812 -3455 5846
rect -3421 5812 -3361 5846
rect -3327 5812 -3311 5846
rect -3135 5812 -3119 5846
rect -3085 5812 -3025 5846
rect -2991 5812 -2975 5846
rect -2799 5812 -2783 5846
rect -2749 5812 -2689 5846
rect -2655 5812 -2639 5846
<< viali >>
rect -4652 8407 -4614 8441
rect -4524 8407 -4486 8441
rect -4248 8407 -4210 8441
rect -4120 8407 -4082 8441
rect -3844 8407 -3806 8441
rect -3716 8407 -3678 8441
rect -3440 8407 -3402 8441
rect -3312 8407 -3274 8441
rect -3036 8407 -2998 8441
rect -2908 8407 -2870 8441
rect -2632 8407 -2594 8441
rect -2504 8407 -2466 8441
rect -4788 8306 -4754 8348
rect -4788 8272 -4754 8306
rect -4788 8238 -4754 8272
rect -4788 8204 -4754 8238
rect -4788 8170 -4754 8204
rect -4788 8136 -4754 8170
rect -4788 8102 -4754 8136
rect -4788 8068 -4754 8102
rect -4788 8034 -4754 8068
rect -4788 8000 -4754 8034
rect -4788 7966 -4754 8000
rect -4788 7932 -4754 7966
rect -4788 7898 -4754 7932
rect -4788 7864 -4754 7898
rect -4788 7830 -4754 7864
rect -4788 7796 -4754 7830
rect -4788 7762 -4754 7796
rect -4788 7728 -4754 7762
rect -4788 7694 -4754 7728
rect -4788 7660 -4754 7694
rect -4788 7626 -4754 7660
rect -4788 7592 -4754 7626
rect -4788 7558 -4754 7592
rect -4788 7524 -4754 7558
rect -4788 7490 -4754 7524
rect -4788 7456 -4754 7490
rect -4788 7422 -4754 7456
rect -4788 7388 -4754 7422
rect -4788 7372 -4754 7388
rect -4714 7372 -4680 8348
rect -4586 7372 -4552 8348
rect -4458 7372 -4424 8348
rect -4384 8332 -4350 8348
rect -4384 8298 -4350 8332
rect -4384 8264 -4350 8298
rect -4384 8230 -4350 8264
rect -4384 8196 -4350 8230
rect -4384 8162 -4350 8196
rect -4384 8128 -4350 8162
rect -4384 8094 -4350 8128
rect -4384 8060 -4350 8094
rect -4384 8026 -4350 8060
rect -4384 7992 -4350 8026
rect -4384 7958 -4350 7992
rect -4384 7924 -4350 7958
rect -4384 7890 -4350 7924
rect -4384 7856 -4350 7890
rect -4384 7822 -4350 7856
rect -4384 7788 -4350 7822
rect -4384 7754 -4350 7788
rect -4384 7720 -4350 7754
rect -4384 7686 -4350 7720
rect -4384 7652 -4350 7686
rect -4384 7618 -4350 7652
rect -4384 7584 -4350 7618
rect -4384 7550 -4350 7584
rect -4384 7516 -4350 7550
rect -4384 7482 -4350 7516
rect -4384 7448 -4350 7482
rect -4384 7414 -4350 7448
rect -4384 7372 -4350 7414
rect -4310 7372 -4276 8348
rect -4182 7372 -4148 8348
rect -4054 7372 -4020 8348
rect -3980 8332 -3946 8348
rect -3980 8298 -3946 8332
rect -3980 8264 -3946 8298
rect -3980 8230 -3946 8264
rect -3980 8196 -3946 8230
rect -3980 8162 -3946 8196
rect -3980 8128 -3946 8162
rect -3980 8094 -3946 8128
rect -3980 8060 -3946 8094
rect -3980 8026 -3946 8060
rect -3980 7992 -3946 8026
rect -3980 7958 -3946 7992
rect -3980 7924 -3946 7958
rect -3980 7890 -3946 7924
rect -3980 7856 -3946 7890
rect -3980 7822 -3946 7856
rect -3980 7788 -3946 7822
rect -3980 7754 -3946 7788
rect -3980 7720 -3946 7754
rect -3980 7686 -3946 7720
rect -3980 7652 -3946 7686
rect -3980 7618 -3946 7652
rect -3980 7584 -3946 7618
rect -3980 7550 -3946 7584
rect -3980 7516 -3946 7550
rect -3980 7482 -3946 7516
rect -3980 7448 -3946 7482
rect -3980 7414 -3946 7448
rect -3980 7372 -3946 7414
rect -3906 7372 -3872 8348
rect -3778 7372 -3744 8348
rect -3650 7372 -3616 8348
rect -3576 8332 -3542 8348
rect -3576 8298 -3542 8332
rect -3576 8264 -3542 8298
rect -3576 8230 -3542 8264
rect -3576 8196 -3542 8230
rect -3576 8162 -3542 8196
rect -3576 8128 -3542 8162
rect -3576 8094 -3542 8128
rect -3576 8060 -3542 8094
rect -3576 8026 -3542 8060
rect -3576 7992 -3542 8026
rect -3576 7958 -3542 7992
rect -3576 7924 -3542 7958
rect -3576 7890 -3542 7924
rect -3576 7856 -3542 7890
rect -3576 7822 -3542 7856
rect -3576 7788 -3542 7822
rect -3576 7754 -3542 7788
rect -3576 7720 -3542 7754
rect -3576 7686 -3542 7720
rect -3576 7652 -3542 7686
rect -3576 7618 -3542 7652
rect -3576 7584 -3542 7618
rect -3576 7550 -3542 7584
rect -3576 7516 -3542 7550
rect -3576 7482 -3542 7516
rect -3576 7448 -3542 7482
rect -3576 7414 -3542 7448
rect -3576 7372 -3542 7414
rect -3502 7372 -3468 8348
rect -3374 7372 -3340 8348
rect -3246 7372 -3212 8348
rect -3172 8332 -3138 8348
rect -3172 8298 -3138 8332
rect -3172 8264 -3138 8298
rect -3172 8230 -3138 8264
rect -3172 8196 -3138 8230
rect -3172 8162 -3138 8196
rect -3172 8128 -3138 8162
rect -3172 8094 -3138 8128
rect -3172 8060 -3138 8094
rect -3172 8026 -3138 8060
rect -3172 7992 -3138 8026
rect -3172 7958 -3138 7992
rect -3172 7924 -3138 7958
rect -3172 7890 -3138 7924
rect -3172 7856 -3138 7890
rect -3172 7822 -3138 7856
rect -3172 7788 -3138 7822
rect -3172 7754 -3138 7788
rect -3172 7720 -3138 7754
rect -3172 7686 -3138 7720
rect -3172 7652 -3138 7686
rect -3172 7618 -3138 7652
rect -3172 7584 -3138 7618
rect -3172 7550 -3138 7584
rect -3172 7516 -3138 7550
rect -3172 7482 -3138 7516
rect -3172 7448 -3138 7482
rect -3172 7414 -3138 7448
rect -3172 7372 -3138 7414
rect -3098 7372 -3064 8348
rect -2970 7372 -2936 8348
rect -2842 7372 -2808 8348
rect -2768 8332 -2734 8348
rect -2768 8298 -2734 8332
rect -2768 8264 -2734 8298
rect -2768 8230 -2734 8264
rect -2768 8196 -2734 8230
rect -2768 8162 -2734 8196
rect -2768 8128 -2734 8162
rect -2768 8094 -2734 8128
rect -2768 8060 -2734 8094
rect -2768 8026 -2734 8060
rect -2768 7992 -2734 8026
rect -2768 7958 -2734 7992
rect -2768 7924 -2734 7958
rect -2768 7890 -2734 7924
rect -2768 7856 -2734 7890
rect -2768 7822 -2734 7856
rect -2768 7788 -2734 7822
rect -2768 7754 -2734 7788
rect -2768 7720 -2734 7754
rect -2768 7686 -2734 7720
rect -2768 7652 -2734 7686
rect -2768 7618 -2734 7652
rect -2768 7584 -2734 7618
rect -2768 7550 -2734 7584
rect -2768 7516 -2734 7550
rect -2768 7482 -2734 7516
rect -2768 7448 -2734 7482
rect -2768 7414 -2734 7448
rect -2768 7372 -2734 7414
rect -2694 7372 -2660 8348
rect -2566 7372 -2532 8348
rect -2438 7372 -2404 8348
rect -2364 8332 -2330 8348
rect -2364 8298 -2330 8332
rect -2364 8264 -2330 8298
rect -2364 8230 -2330 8264
rect -2364 8196 -2330 8230
rect -2364 8162 -2330 8196
rect -2364 8128 -2330 8162
rect -2364 8094 -2330 8128
rect -2364 8060 -2330 8094
rect -2364 8026 -2330 8060
rect -2364 7992 -2330 8026
rect -2364 7958 -2330 7992
rect -2364 7924 -2330 7958
rect -2364 7890 -2330 7924
rect -2364 7856 -2330 7890
rect -2364 7822 -2330 7856
rect -2364 7788 -2330 7822
rect -2364 7754 -2330 7788
rect -2364 7720 -2330 7754
rect -2364 7686 -2330 7720
rect -2364 7652 -2330 7686
rect -2364 7618 -2330 7652
rect -2364 7584 -2330 7618
rect -2364 7550 -2330 7584
rect -2364 7516 -2330 7550
rect -2364 7482 -2330 7516
rect -2364 7448 -2330 7482
rect -2364 7414 -2330 7448
rect -2364 7372 -2330 7414
rect 610 8356 644 8398
rect 610 8322 644 8356
rect 610 8288 644 8322
rect 610 8254 644 8288
rect 610 8220 644 8254
rect 610 8186 644 8220
rect 610 8152 644 8186
rect 610 8118 644 8152
rect 610 8084 644 8118
rect 610 8050 644 8084
rect 610 8016 644 8050
rect 610 7982 644 8016
rect 610 7948 644 7982
rect 610 7914 644 7948
rect 610 7880 644 7914
rect 610 7846 644 7880
rect 610 7812 644 7846
rect 610 7778 644 7812
rect 610 7744 644 7778
rect 610 7710 644 7744
rect 610 7676 644 7710
rect 610 7642 644 7676
rect 610 7608 644 7642
rect 610 7574 644 7608
rect 610 7540 644 7574
rect 610 7506 644 7540
rect 610 7472 644 7506
rect 610 7438 644 7472
rect 610 7422 644 7438
rect 684 7422 718 8398
rect 812 7422 846 8398
rect 940 7422 974 8398
rect 1014 8382 1048 8398
rect 1014 8348 1048 8382
rect 1014 8314 1048 8348
rect 1014 8280 1048 8314
rect 1014 8246 1048 8280
rect 1014 8212 1048 8246
rect 1014 8178 1048 8212
rect 1014 8144 1048 8178
rect 1014 8110 1048 8144
rect 1014 8076 1048 8110
rect 1014 8042 1048 8076
rect 1014 8008 1048 8042
rect 1014 7974 1048 8008
rect 1014 7940 1048 7974
rect 1014 7906 1048 7940
rect 1014 7872 1048 7906
rect 1014 7838 1048 7872
rect 1014 7804 1048 7838
rect 1014 7770 1048 7804
rect 1014 7736 1048 7770
rect 1014 7702 1048 7736
rect 1014 7668 1048 7702
rect 1014 7634 1048 7668
rect 1014 7600 1048 7634
rect 1014 7566 1048 7600
rect 1014 7532 1048 7566
rect 1014 7498 1048 7532
rect 1014 7464 1048 7498
rect 1014 7422 1048 7464
rect 1088 7422 1122 8398
rect 1216 7422 1250 8398
rect 1344 7422 1378 8398
rect 1418 8382 1452 8398
rect 1418 8348 1452 8382
rect 1418 8314 1452 8348
rect 1418 8280 1452 8314
rect 1418 8246 1452 8280
rect 1418 8212 1452 8246
rect 1418 8178 1452 8212
rect 1418 8144 1452 8178
rect 1418 8110 1452 8144
rect 1418 8076 1452 8110
rect 1418 8042 1452 8076
rect 1418 8008 1452 8042
rect 1418 7974 1452 8008
rect 1418 7940 1452 7974
rect 1418 7906 1452 7940
rect 1418 7872 1452 7906
rect 1418 7838 1452 7872
rect 1418 7804 1452 7838
rect 1418 7770 1452 7804
rect 1418 7736 1452 7770
rect 1418 7702 1452 7736
rect 1418 7668 1452 7702
rect 1418 7634 1452 7668
rect 1418 7600 1452 7634
rect 1418 7566 1452 7600
rect 1418 7532 1452 7566
rect 1418 7498 1452 7532
rect 1418 7464 1452 7498
rect 1418 7422 1452 7464
rect 1492 7422 1526 8398
rect 1620 7422 1654 8398
rect 1748 7422 1782 8398
rect 1822 8382 1856 8398
rect 1822 8348 1856 8382
rect 1822 8314 1856 8348
rect 1822 8280 1856 8314
rect 1822 8246 1856 8280
rect 1822 8212 1856 8246
rect 1822 8178 1856 8212
rect 1822 8144 1856 8178
rect 1822 8110 1856 8144
rect 1822 8076 1856 8110
rect 1822 8042 1856 8076
rect 1822 8008 1856 8042
rect 1822 7974 1856 8008
rect 1822 7940 1856 7974
rect 1822 7906 1856 7940
rect 1822 7872 1856 7906
rect 1822 7838 1856 7872
rect 1822 7804 1856 7838
rect 1822 7770 1856 7804
rect 1822 7736 1856 7770
rect 1822 7702 1856 7736
rect 1822 7668 1856 7702
rect 1822 7634 1856 7668
rect 1822 7600 1856 7634
rect 1822 7566 1856 7600
rect 1822 7532 1856 7566
rect 1822 7498 1856 7532
rect 1822 7464 1856 7498
rect 1822 7422 1856 7464
rect 1896 7422 1930 8398
rect 2024 7422 2058 8398
rect 2152 7422 2186 8398
rect 2226 8382 2260 8398
rect 2226 8348 2260 8382
rect 2226 8314 2260 8348
rect 2226 8280 2260 8314
rect 2226 8246 2260 8280
rect 2226 8212 2260 8246
rect 2226 8178 2260 8212
rect 2226 8144 2260 8178
rect 2226 8110 2260 8144
rect 2226 8076 2260 8110
rect 2226 8042 2260 8076
rect 2226 8008 2260 8042
rect 2226 7974 2260 8008
rect 2226 7940 2260 7974
rect 2226 7906 2260 7940
rect 2226 7872 2260 7906
rect 2226 7838 2260 7872
rect 2226 7804 2260 7838
rect 2226 7770 2260 7804
rect 2226 7736 2260 7770
rect 2226 7702 2260 7736
rect 2226 7668 2260 7702
rect 2226 7634 2260 7668
rect 2226 7600 2260 7634
rect 2226 7566 2260 7600
rect 2226 7532 2260 7566
rect 2226 7498 2260 7532
rect 2226 7464 2260 7498
rect 2226 7422 2260 7464
rect 2300 7422 2334 8398
rect 2428 7422 2462 8398
rect 2556 7422 2590 8398
rect 2630 8382 2664 8398
rect 2630 8348 2664 8382
rect 2630 8314 2664 8348
rect 2630 8280 2664 8314
rect 2630 8246 2664 8280
rect 2630 8212 2664 8246
rect 2630 8178 2664 8212
rect 2630 8144 2664 8178
rect 2630 8110 2664 8144
rect 2630 8076 2664 8110
rect 2630 8042 2664 8076
rect 2630 8008 2664 8042
rect 2630 7974 2664 8008
rect 2630 7940 2664 7974
rect 2630 7906 2664 7940
rect 2630 7872 2664 7906
rect 2630 7838 2664 7872
rect 2630 7804 2664 7838
rect 2630 7770 2664 7804
rect 2630 7736 2664 7770
rect 2630 7702 2664 7736
rect 2630 7668 2664 7702
rect 2630 7634 2664 7668
rect 2630 7600 2664 7634
rect 2630 7566 2664 7600
rect 2630 7532 2664 7566
rect 2630 7498 2664 7532
rect 2630 7464 2664 7498
rect 2630 7422 2664 7464
rect 2704 7422 2738 8398
rect 2832 7422 2866 8398
rect 2960 7422 2994 8398
rect 3034 8382 3068 8398
rect 3034 8348 3068 8382
rect 3034 8314 3068 8348
rect 3034 8280 3068 8314
rect 3034 8246 3068 8280
rect 3034 8212 3068 8246
rect 3034 8178 3068 8212
rect 3034 8144 3068 8178
rect 3034 8110 3068 8144
rect 3034 8076 3068 8110
rect 3034 8042 3068 8076
rect 3034 8008 3068 8042
rect 3034 7974 3068 8008
rect 3034 7940 3068 7974
rect 3034 7906 3068 7940
rect 3034 7872 3068 7906
rect 3034 7838 3068 7872
rect 3034 7804 3068 7838
rect 3034 7770 3068 7804
rect 3034 7736 3068 7770
rect 3034 7702 3068 7736
rect 3034 7668 3068 7702
rect 3034 7634 3068 7668
rect 3034 7600 3068 7634
rect 3034 7566 3068 7600
rect 3034 7532 3068 7566
rect 3034 7498 3068 7532
rect 3034 7464 3068 7498
rect 3034 7422 3068 7464
rect 6980 8356 7014 8398
rect 6980 8322 7014 8356
rect 6980 8288 7014 8322
rect 6980 8254 7014 8288
rect 6980 8220 7014 8254
rect 6980 8186 7014 8220
rect 6980 8152 7014 8186
rect 6980 8118 7014 8152
rect 6980 8084 7014 8118
rect 6980 8050 7014 8084
rect 6980 8016 7014 8050
rect 6980 7982 7014 8016
rect 6980 7948 7014 7982
rect 6980 7914 7014 7948
rect 6980 7880 7014 7914
rect 6980 7846 7014 7880
rect 6980 7812 7014 7846
rect 6980 7778 7014 7812
rect 6980 7744 7014 7778
rect 6980 7710 7014 7744
rect 6980 7676 7014 7710
rect 6980 7642 7014 7676
rect 6980 7608 7014 7642
rect 6980 7574 7014 7608
rect 6980 7540 7014 7574
rect 6980 7506 7014 7540
rect 6980 7472 7014 7506
rect 6980 7438 7014 7472
rect 6980 7422 7014 7438
rect 7054 7422 7088 8398
rect 7182 7422 7216 8398
rect 7310 7422 7344 8398
rect 7384 8382 7418 8398
rect 7384 8348 7418 8382
rect 7384 8314 7418 8348
rect 7384 8280 7418 8314
rect 7384 8246 7418 8280
rect 7384 8212 7418 8246
rect 7384 8178 7418 8212
rect 7384 8144 7418 8178
rect 7384 8110 7418 8144
rect 7384 8076 7418 8110
rect 7384 8042 7418 8076
rect 7384 8008 7418 8042
rect 7384 7974 7418 8008
rect 7384 7940 7418 7974
rect 7384 7906 7418 7940
rect 7384 7872 7418 7906
rect 7384 7838 7418 7872
rect 7384 7804 7418 7838
rect 7384 7770 7418 7804
rect 7384 7736 7418 7770
rect 7384 7702 7418 7736
rect 7384 7668 7418 7702
rect 7384 7634 7418 7668
rect 7384 7600 7418 7634
rect 7384 7566 7418 7600
rect 7384 7532 7418 7566
rect 7384 7498 7418 7532
rect 7384 7464 7418 7498
rect 7384 7422 7418 7464
rect 7458 7422 7492 8398
rect 7586 7422 7620 8398
rect 7714 7422 7748 8398
rect 7788 8382 7822 8398
rect 7788 8348 7822 8382
rect 7788 8314 7822 8348
rect 7788 8280 7822 8314
rect 7788 8246 7822 8280
rect 7788 8212 7822 8246
rect 7788 8178 7822 8212
rect 7788 8144 7822 8178
rect 7788 8110 7822 8144
rect 7788 8076 7822 8110
rect 7788 8042 7822 8076
rect 7788 8008 7822 8042
rect 7788 7974 7822 8008
rect 7788 7940 7822 7974
rect 7788 7906 7822 7940
rect 7788 7872 7822 7906
rect 7788 7838 7822 7872
rect 7788 7804 7822 7838
rect 7788 7770 7822 7804
rect 7788 7736 7822 7770
rect 7788 7702 7822 7736
rect 7788 7668 7822 7702
rect 7788 7634 7822 7668
rect 7788 7600 7822 7634
rect 7788 7566 7822 7600
rect 7788 7532 7822 7566
rect 7788 7498 7822 7532
rect 7788 7464 7822 7498
rect 7788 7422 7822 7464
rect 7862 7422 7896 8398
rect 7990 7422 8024 8398
rect 8118 7422 8152 8398
rect 8192 8382 8226 8398
rect 8192 8348 8226 8382
rect 8192 8314 8226 8348
rect 8192 8280 8226 8314
rect 8192 8246 8226 8280
rect 8192 8212 8226 8246
rect 8192 8178 8226 8212
rect 8192 8144 8226 8178
rect 8192 8110 8226 8144
rect 8192 8076 8226 8110
rect 8192 8042 8226 8076
rect 8192 8008 8226 8042
rect 8192 7974 8226 8008
rect 8192 7940 8226 7974
rect 8192 7906 8226 7940
rect 8192 7872 8226 7906
rect 8192 7838 8226 7872
rect 8192 7804 8226 7838
rect 8192 7770 8226 7804
rect 8192 7736 8226 7770
rect 8192 7702 8226 7736
rect 8192 7668 8226 7702
rect 8192 7634 8226 7668
rect 8192 7600 8226 7634
rect 8192 7566 8226 7600
rect 8192 7532 8226 7566
rect 8192 7498 8226 7532
rect 8192 7464 8226 7498
rect 8192 7422 8226 7464
rect 8266 7422 8300 8398
rect 8394 7422 8428 8398
rect 8522 7422 8556 8398
rect 8596 8382 8630 8398
rect 8596 8348 8630 8382
rect 8596 8314 8630 8348
rect 8596 8280 8630 8314
rect 8596 8246 8630 8280
rect 8596 8212 8630 8246
rect 8596 8178 8630 8212
rect 8596 8144 8630 8178
rect 8596 8110 8630 8144
rect 8596 8076 8630 8110
rect 8596 8042 8630 8076
rect 8596 8008 8630 8042
rect 8596 7974 8630 8008
rect 8596 7940 8630 7974
rect 8596 7906 8630 7940
rect 8596 7872 8630 7906
rect 8596 7838 8630 7872
rect 8596 7804 8630 7838
rect 8596 7770 8630 7804
rect 8596 7736 8630 7770
rect 8596 7702 8630 7736
rect 8596 7668 8630 7702
rect 8596 7634 8630 7668
rect 8596 7600 8630 7634
rect 8596 7566 8630 7600
rect 8596 7532 8630 7566
rect 8596 7498 8630 7532
rect 8596 7464 8630 7498
rect 8596 7422 8630 7464
rect 8670 7422 8704 8398
rect 8798 7422 8832 8398
rect 8926 7422 8960 8398
rect 9000 8382 9034 8398
rect 9000 8348 9034 8382
rect 9000 8314 9034 8348
rect 9000 8280 9034 8314
rect 9000 8246 9034 8280
rect 9000 8212 9034 8246
rect 9000 8178 9034 8212
rect 9000 8144 9034 8178
rect 9000 8110 9034 8144
rect 9000 8076 9034 8110
rect 9000 8042 9034 8076
rect 9000 8008 9034 8042
rect 9000 7974 9034 8008
rect 9000 7940 9034 7974
rect 9000 7906 9034 7940
rect 9000 7872 9034 7906
rect 9000 7838 9034 7872
rect 9000 7804 9034 7838
rect 9000 7770 9034 7804
rect 9000 7736 9034 7770
rect 9000 7702 9034 7736
rect 9000 7668 9034 7702
rect 9000 7634 9034 7668
rect 9000 7600 9034 7634
rect 9000 7566 9034 7600
rect 9000 7532 9034 7566
rect 9000 7498 9034 7532
rect 9000 7464 9034 7498
rect 9000 7422 9034 7464
rect 9074 7422 9108 8398
rect 9202 7422 9236 8398
rect 9330 7422 9364 8398
rect 9404 8382 9438 8398
rect 9404 8348 9438 8382
rect 9404 8314 9438 8348
rect 9404 8280 9438 8314
rect 9404 8246 9438 8280
rect 9404 8212 9438 8246
rect 9404 8178 9438 8212
rect 9404 8144 9438 8178
rect 9404 8110 9438 8144
rect 9404 8076 9438 8110
rect 9404 8042 9438 8076
rect 9404 8008 9438 8042
rect 9404 7974 9438 8008
rect 9404 7940 9438 7974
rect 9404 7906 9438 7940
rect 9404 7872 9438 7906
rect 9404 7838 9438 7872
rect 9404 7804 9438 7838
rect 9404 7770 9438 7804
rect 9404 7736 9438 7770
rect 9404 7702 9438 7736
rect 9404 7668 9438 7702
rect 9404 7634 9438 7668
rect 9404 7600 9438 7634
rect 9404 7566 9438 7600
rect 9404 7532 9438 7566
rect 9404 7498 9438 7532
rect 9404 7464 9438 7498
rect 9404 7422 9438 7464
rect 13350 8356 13384 8398
rect 13350 8322 13384 8356
rect 13350 8288 13384 8322
rect 13350 8254 13384 8288
rect 13350 8220 13384 8254
rect 13350 8186 13384 8220
rect 13350 8152 13384 8186
rect 13350 8118 13384 8152
rect 13350 8084 13384 8118
rect 13350 8050 13384 8084
rect 13350 8016 13384 8050
rect 13350 7982 13384 8016
rect 13350 7948 13384 7982
rect 13350 7914 13384 7948
rect 13350 7880 13384 7914
rect 13350 7846 13384 7880
rect 13350 7812 13384 7846
rect 13350 7778 13384 7812
rect 13350 7744 13384 7778
rect 13350 7710 13384 7744
rect 13350 7676 13384 7710
rect 13350 7642 13384 7676
rect 13350 7608 13384 7642
rect 13350 7574 13384 7608
rect 13350 7540 13384 7574
rect 13350 7506 13384 7540
rect 13350 7472 13384 7506
rect 13350 7438 13384 7472
rect 13350 7422 13384 7438
rect 13424 7422 13458 8398
rect 13552 7422 13586 8398
rect 13680 7422 13714 8398
rect 13754 8382 13788 8398
rect 13754 8348 13788 8382
rect 13754 8314 13788 8348
rect 13754 8280 13788 8314
rect 13754 8246 13788 8280
rect 13754 8212 13788 8246
rect 13754 8178 13788 8212
rect 13754 8144 13788 8178
rect 13754 8110 13788 8144
rect 13754 8076 13788 8110
rect 13754 8042 13788 8076
rect 13754 8008 13788 8042
rect 13754 7974 13788 8008
rect 13754 7940 13788 7974
rect 13754 7906 13788 7940
rect 13754 7872 13788 7906
rect 13754 7838 13788 7872
rect 13754 7804 13788 7838
rect 13754 7770 13788 7804
rect 13754 7736 13788 7770
rect 13754 7702 13788 7736
rect 13754 7668 13788 7702
rect 13754 7634 13788 7668
rect 13754 7600 13788 7634
rect 13754 7566 13788 7600
rect 13754 7532 13788 7566
rect 13754 7498 13788 7532
rect 13754 7464 13788 7498
rect 13754 7422 13788 7464
rect 13828 7422 13862 8398
rect 13956 7422 13990 8398
rect 14084 7422 14118 8398
rect 14158 8382 14192 8398
rect 14158 8348 14192 8382
rect 14158 8314 14192 8348
rect 14158 8280 14192 8314
rect 14158 8246 14192 8280
rect 14158 8212 14192 8246
rect 14158 8178 14192 8212
rect 14158 8144 14192 8178
rect 14158 8110 14192 8144
rect 14158 8076 14192 8110
rect 14158 8042 14192 8076
rect 14158 8008 14192 8042
rect 14158 7974 14192 8008
rect 14158 7940 14192 7974
rect 14158 7906 14192 7940
rect 14158 7872 14192 7906
rect 14158 7838 14192 7872
rect 14158 7804 14192 7838
rect 14158 7770 14192 7804
rect 14158 7736 14192 7770
rect 14158 7702 14192 7736
rect 14158 7668 14192 7702
rect 14158 7634 14192 7668
rect 14158 7600 14192 7634
rect 14158 7566 14192 7600
rect 14158 7532 14192 7566
rect 14158 7498 14192 7532
rect 14158 7464 14192 7498
rect 14158 7422 14192 7464
rect 14232 7422 14266 8398
rect 14360 7422 14394 8398
rect 14488 7422 14522 8398
rect 14562 8382 14596 8398
rect 14562 8348 14596 8382
rect 14562 8314 14596 8348
rect 14562 8280 14596 8314
rect 14562 8246 14596 8280
rect 14562 8212 14596 8246
rect 14562 8178 14596 8212
rect 14562 8144 14596 8178
rect 14562 8110 14596 8144
rect 14562 8076 14596 8110
rect 14562 8042 14596 8076
rect 14562 8008 14596 8042
rect 14562 7974 14596 8008
rect 14562 7940 14596 7974
rect 14562 7906 14596 7940
rect 14562 7872 14596 7906
rect 14562 7838 14596 7872
rect 14562 7804 14596 7838
rect 14562 7770 14596 7804
rect 14562 7736 14596 7770
rect 14562 7702 14596 7736
rect 14562 7668 14596 7702
rect 14562 7634 14596 7668
rect 14562 7600 14596 7634
rect 14562 7566 14596 7600
rect 14562 7532 14596 7566
rect 14562 7498 14596 7532
rect 14562 7464 14596 7498
rect 14562 7422 14596 7464
rect 14636 7422 14670 8398
rect 14764 7422 14798 8398
rect 14892 7422 14926 8398
rect 14966 8382 15000 8398
rect 14966 8348 15000 8382
rect 14966 8314 15000 8348
rect 14966 8280 15000 8314
rect 14966 8246 15000 8280
rect 14966 8212 15000 8246
rect 14966 8178 15000 8212
rect 14966 8144 15000 8178
rect 14966 8110 15000 8144
rect 14966 8076 15000 8110
rect 14966 8042 15000 8076
rect 14966 8008 15000 8042
rect 14966 7974 15000 8008
rect 14966 7940 15000 7974
rect 14966 7906 15000 7940
rect 14966 7872 15000 7906
rect 14966 7838 15000 7872
rect 14966 7804 15000 7838
rect 14966 7770 15000 7804
rect 14966 7736 15000 7770
rect 14966 7702 15000 7736
rect 14966 7668 15000 7702
rect 14966 7634 15000 7668
rect 14966 7600 15000 7634
rect 14966 7566 15000 7600
rect 14966 7532 15000 7566
rect 14966 7498 15000 7532
rect 14966 7464 15000 7498
rect 14966 7422 15000 7464
rect 15040 7422 15074 8398
rect 15168 7422 15202 8398
rect 15296 7422 15330 8398
rect 15370 8382 15404 8398
rect 15370 8348 15404 8382
rect 15370 8314 15404 8348
rect 15370 8280 15404 8314
rect 15370 8246 15404 8280
rect 15370 8212 15404 8246
rect 15370 8178 15404 8212
rect 15370 8144 15404 8178
rect 15370 8110 15404 8144
rect 15370 8076 15404 8110
rect 15370 8042 15404 8076
rect 15370 8008 15404 8042
rect 15370 7974 15404 8008
rect 15370 7940 15404 7974
rect 15370 7906 15404 7940
rect 15370 7872 15404 7906
rect 15370 7838 15404 7872
rect 15370 7804 15404 7838
rect 15370 7770 15404 7804
rect 15370 7736 15404 7770
rect 15370 7702 15404 7736
rect 15370 7668 15404 7702
rect 15370 7634 15404 7668
rect 15370 7600 15404 7634
rect 15370 7566 15404 7600
rect 15370 7532 15404 7566
rect 15370 7498 15404 7532
rect 15370 7464 15404 7498
rect 15370 7422 15404 7464
rect 15444 7422 15478 8398
rect 15572 7422 15606 8398
rect 15700 7422 15734 8398
rect 15774 8382 15808 8398
rect 15774 8348 15808 8382
rect 15774 8314 15808 8348
rect 15774 8280 15808 8314
rect 15774 8246 15808 8280
rect 15774 8212 15808 8246
rect 15774 8178 15808 8212
rect 15774 8144 15808 8178
rect 15774 8110 15808 8144
rect 15774 8076 15808 8110
rect 15774 8042 15808 8076
rect 15774 8008 15808 8042
rect 15774 7974 15808 8008
rect 15774 7940 15808 7974
rect 15774 7906 15808 7940
rect 15774 7872 15808 7906
rect 15774 7838 15808 7872
rect 15774 7804 15808 7838
rect 15774 7770 15808 7804
rect 15774 7736 15808 7770
rect 15774 7702 15808 7736
rect 15774 7668 15808 7702
rect 15774 7634 15808 7668
rect 15774 7600 15808 7634
rect 15774 7566 15808 7600
rect 15774 7532 15808 7566
rect 15774 7498 15808 7532
rect 15774 7464 15808 7498
rect 15774 7422 15808 7464
rect 19720 8356 19754 8398
rect 19720 8322 19754 8356
rect 19720 8288 19754 8322
rect 19720 8254 19754 8288
rect 19720 8220 19754 8254
rect 19720 8186 19754 8220
rect 19720 8152 19754 8186
rect 19720 8118 19754 8152
rect 19720 8084 19754 8118
rect 19720 8050 19754 8084
rect 19720 8016 19754 8050
rect 19720 7982 19754 8016
rect 19720 7948 19754 7982
rect 19720 7914 19754 7948
rect 19720 7880 19754 7914
rect 19720 7846 19754 7880
rect 19720 7812 19754 7846
rect 19720 7778 19754 7812
rect 19720 7744 19754 7778
rect 19720 7710 19754 7744
rect 19720 7676 19754 7710
rect 19720 7642 19754 7676
rect 19720 7608 19754 7642
rect 19720 7574 19754 7608
rect 19720 7540 19754 7574
rect 19720 7506 19754 7540
rect 19720 7472 19754 7506
rect 19720 7438 19754 7472
rect 19720 7422 19754 7438
rect 19794 7422 19828 8398
rect 19922 7422 19956 8398
rect 20050 7422 20084 8398
rect 20124 8382 20158 8398
rect 20124 8348 20158 8382
rect 20124 8314 20158 8348
rect 20124 8280 20158 8314
rect 20124 8246 20158 8280
rect 20124 8212 20158 8246
rect 20124 8178 20158 8212
rect 20124 8144 20158 8178
rect 20124 8110 20158 8144
rect 20124 8076 20158 8110
rect 20124 8042 20158 8076
rect 20124 8008 20158 8042
rect 20124 7974 20158 8008
rect 20124 7940 20158 7974
rect 20124 7906 20158 7940
rect 20124 7872 20158 7906
rect 20124 7838 20158 7872
rect 20124 7804 20158 7838
rect 20124 7770 20158 7804
rect 20124 7736 20158 7770
rect 20124 7702 20158 7736
rect 20124 7668 20158 7702
rect 20124 7634 20158 7668
rect 20124 7600 20158 7634
rect 20124 7566 20158 7600
rect 20124 7532 20158 7566
rect 20124 7498 20158 7532
rect 20124 7464 20158 7498
rect 20124 7422 20158 7464
rect 20198 7422 20232 8398
rect 20326 7422 20360 8398
rect 20454 7422 20488 8398
rect 20528 8382 20562 8398
rect 20528 8348 20562 8382
rect 20528 8314 20562 8348
rect 20528 8280 20562 8314
rect 20528 8246 20562 8280
rect 20528 8212 20562 8246
rect 20528 8178 20562 8212
rect 20528 8144 20562 8178
rect 20528 8110 20562 8144
rect 20528 8076 20562 8110
rect 20528 8042 20562 8076
rect 20528 8008 20562 8042
rect 20528 7974 20562 8008
rect 20528 7940 20562 7974
rect 20528 7906 20562 7940
rect 20528 7872 20562 7906
rect 20528 7838 20562 7872
rect 20528 7804 20562 7838
rect 20528 7770 20562 7804
rect 20528 7736 20562 7770
rect 20528 7702 20562 7736
rect 20528 7668 20562 7702
rect 20528 7634 20562 7668
rect 20528 7600 20562 7634
rect 20528 7566 20562 7600
rect 20528 7532 20562 7566
rect 20528 7498 20562 7532
rect 20528 7464 20562 7498
rect 20528 7422 20562 7464
rect 20602 7422 20636 8398
rect 20730 7422 20764 8398
rect 20858 7422 20892 8398
rect 20932 8382 20966 8398
rect 20932 8348 20966 8382
rect 20932 8314 20966 8348
rect 20932 8280 20966 8314
rect 20932 8246 20966 8280
rect 20932 8212 20966 8246
rect 20932 8178 20966 8212
rect 20932 8144 20966 8178
rect 20932 8110 20966 8144
rect 20932 8076 20966 8110
rect 20932 8042 20966 8076
rect 20932 8008 20966 8042
rect 20932 7974 20966 8008
rect 20932 7940 20966 7974
rect 20932 7906 20966 7940
rect 20932 7872 20966 7906
rect 20932 7838 20966 7872
rect 20932 7804 20966 7838
rect 20932 7770 20966 7804
rect 20932 7736 20966 7770
rect 20932 7702 20966 7736
rect 20932 7668 20966 7702
rect 20932 7634 20966 7668
rect 20932 7600 20966 7634
rect 20932 7566 20966 7600
rect 20932 7532 20966 7566
rect 20932 7498 20966 7532
rect 20932 7464 20966 7498
rect 20932 7422 20966 7464
rect 21006 7422 21040 8398
rect 21134 7422 21168 8398
rect 21262 7422 21296 8398
rect 21336 8382 21370 8398
rect 21336 8348 21370 8382
rect 21336 8314 21370 8348
rect 21336 8280 21370 8314
rect 21336 8246 21370 8280
rect 21336 8212 21370 8246
rect 21336 8178 21370 8212
rect 21336 8144 21370 8178
rect 21336 8110 21370 8144
rect 21336 8076 21370 8110
rect 21336 8042 21370 8076
rect 21336 8008 21370 8042
rect 21336 7974 21370 8008
rect 21336 7940 21370 7974
rect 21336 7906 21370 7940
rect 21336 7872 21370 7906
rect 21336 7838 21370 7872
rect 21336 7804 21370 7838
rect 21336 7770 21370 7804
rect 21336 7736 21370 7770
rect 21336 7702 21370 7736
rect 21336 7668 21370 7702
rect 21336 7634 21370 7668
rect 21336 7600 21370 7634
rect 21336 7566 21370 7600
rect 21336 7532 21370 7566
rect 21336 7498 21370 7532
rect 21336 7464 21370 7498
rect 21336 7422 21370 7464
rect 21410 7422 21444 8398
rect 21538 7422 21572 8398
rect 21666 7422 21700 8398
rect 21740 8382 21774 8398
rect 21740 8348 21774 8382
rect 21740 8314 21774 8348
rect 21740 8280 21774 8314
rect 21740 8246 21774 8280
rect 21740 8212 21774 8246
rect 21740 8178 21774 8212
rect 21740 8144 21774 8178
rect 21740 8110 21774 8144
rect 21740 8076 21774 8110
rect 21740 8042 21774 8076
rect 21740 8008 21774 8042
rect 21740 7974 21774 8008
rect 21740 7940 21774 7974
rect 21740 7906 21774 7940
rect 21740 7872 21774 7906
rect 21740 7838 21774 7872
rect 21740 7804 21774 7838
rect 21740 7770 21774 7804
rect 21740 7736 21774 7770
rect 21740 7702 21774 7736
rect 21740 7668 21774 7702
rect 21740 7634 21774 7668
rect 21740 7600 21774 7634
rect 21740 7566 21774 7600
rect 21740 7532 21774 7566
rect 21740 7498 21774 7532
rect 21740 7464 21774 7498
rect 21740 7422 21774 7464
rect 21814 7422 21848 8398
rect 21942 7422 21976 8398
rect 22070 7422 22104 8398
rect 22144 8382 22178 8398
rect 22144 8348 22178 8382
rect 22144 8314 22178 8348
rect 22144 8280 22178 8314
rect 22144 8246 22178 8280
rect 22144 8212 22178 8246
rect 22144 8178 22178 8212
rect 22144 8144 22178 8178
rect 22144 8110 22178 8144
rect 22144 8076 22178 8110
rect 22144 8042 22178 8076
rect 22144 8008 22178 8042
rect 22144 7974 22178 8008
rect 22144 7940 22178 7974
rect 22144 7906 22178 7940
rect 22144 7872 22178 7906
rect 22144 7838 22178 7872
rect 22144 7804 22178 7838
rect 22144 7770 22178 7804
rect 22144 7736 22178 7770
rect 22144 7702 22178 7736
rect 22144 7668 22178 7702
rect 22144 7634 22178 7668
rect 22144 7600 22178 7634
rect 22144 7566 22178 7600
rect 22144 7532 22178 7566
rect 22144 7498 22178 7532
rect 22144 7464 22178 7498
rect 22144 7422 22178 7464
rect 28978 8356 29012 8398
rect 28978 8322 29012 8356
rect 28978 8288 29012 8322
rect 28978 8254 29012 8288
rect 28978 8220 29012 8254
rect 28978 8186 29012 8220
rect 28978 8152 29012 8186
rect 28978 8118 29012 8152
rect 28978 8084 29012 8118
rect 28978 8050 29012 8084
rect 28978 8016 29012 8050
rect 28978 7982 29012 8016
rect 28978 7948 29012 7982
rect 28978 7914 29012 7948
rect 28978 7880 29012 7914
rect 28978 7846 29012 7880
rect 28978 7812 29012 7846
rect 28978 7778 29012 7812
rect 28978 7744 29012 7778
rect 28978 7710 29012 7744
rect 28978 7676 29012 7710
rect 28978 7642 29012 7676
rect 28978 7608 29012 7642
rect 28978 7574 29012 7608
rect 28978 7540 29012 7574
rect 28978 7506 29012 7540
rect 28978 7472 29012 7506
rect 28978 7438 29012 7472
rect 28978 7422 29012 7438
rect 29052 7422 29086 8398
rect 29180 7422 29214 8398
rect 29308 7422 29342 8398
rect 29382 8382 29416 8398
rect 29382 8348 29416 8382
rect 29382 8314 29416 8348
rect 29382 8280 29416 8314
rect 29382 8246 29416 8280
rect 29382 8212 29416 8246
rect 29382 8178 29416 8212
rect 29382 8144 29416 8178
rect 29382 8110 29416 8144
rect 29382 8076 29416 8110
rect 29382 8042 29416 8076
rect 29382 8008 29416 8042
rect 29382 7974 29416 8008
rect 29382 7940 29416 7974
rect 29382 7906 29416 7940
rect 29382 7872 29416 7906
rect 29382 7838 29416 7872
rect 29382 7804 29416 7838
rect 29382 7770 29416 7804
rect 29382 7736 29416 7770
rect 29382 7702 29416 7736
rect 29382 7668 29416 7702
rect 29382 7634 29416 7668
rect 29382 7600 29416 7634
rect 29382 7566 29416 7600
rect 29382 7532 29416 7566
rect 29382 7498 29416 7532
rect 29382 7464 29416 7498
rect 29382 7422 29416 7464
rect 29456 7422 29490 8398
rect 29584 7422 29618 8398
rect 29712 7422 29746 8398
rect 29786 8382 29820 8398
rect 29786 8348 29820 8382
rect 29786 8314 29820 8348
rect 29786 8280 29820 8314
rect 29786 8246 29820 8280
rect 29786 8212 29820 8246
rect 29786 8178 29820 8212
rect 29786 8144 29820 8178
rect 29786 8110 29820 8144
rect 29786 8076 29820 8110
rect 29786 8042 29820 8076
rect 29786 8008 29820 8042
rect 29786 7974 29820 8008
rect 29786 7940 29820 7974
rect 29786 7906 29820 7940
rect 29786 7872 29820 7906
rect 29786 7838 29820 7872
rect 29786 7804 29820 7838
rect 29786 7770 29820 7804
rect 29786 7736 29820 7770
rect 29786 7702 29820 7736
rect 29786 7668 29820 7702
rect 29786 7634 29820 7668
rect 29786 7600 29820 7634
rect 29786 7566 29820 7600
rect 29786 7532 29820 7566
rect 29786 7498 29820 7532
rect 29786 7464 29820 7498
rect 29786 7422 29820 7464
rect 29860 7422 29894 8398
rect 29988 7422 30022 8398
rect 30116 7422 30150 8398
rect 30190 8382 30224 8398
rect 30190 8348 30224 8382
rect 30190 8314 30224 8348
rect 30190 8280 30224 8314
rect 30190 8246 30224 8280
rect 30190 8212 30224 8246
rect 30190 8178 30224 8212
rect 30190 8144 30224 8178
rect 30190 8110 30224 8144
rect 30190 8076 30224 8110
rect 30190 8042 30224 8076
rect 30190 8008 30224 8042
rect 30190 7974 30224 8008
rect 30190 7940 30224 7974
rect 30190 7906 30224 7940
rect 30190 7872 30224 7906
rect 30190 7838 30224 7872
rect 30190 7804 30224 7838
rect 30190 7770 30224 7804
rect 30190 7736 30224 7770
rect 30190 7702 30224 7736
rect 30190 7668 30224 7702
rect 30190 7634 30224 7668
rect 30190 7600 30224 7634
rect 30190 7566 30224 7600
rect 30190 7532 30224 7566
rect 30190 7498 30224 7532
rect 30190 7464 30224 7498
rect 30190 7422 30224 7464
rect 30264 7422 30298 8398
rect 30392 7422 30426 8398
rect 30520 7422 30554 8398
rect 30594 8382 30628 8398
rect 30594 8348 30628 8382
rect 30594 8314 30628 8348
rect 30594 8280 30628 8314
rect 30594 8246 30628 8280
rect 30594 8212 30628 8246
rect 30594 8178 30628 8212
rect 30594 8144 30628 8178
rect 30594 8110 30628 8144
rect 30594 8076 30628 8110
rect 30594 8042 30628 8076
rect 30594 8008 30628 8042
rect 30594 7974 30628 8008
rect 30594 7940 30628 7974
rect 30594 7906 30628 7940
rect 30594 7872 30628 7906
rect 30594 7838 30628 7872
rect 30594 7804 30628 7838
rect 30594 7770 30628 7804
rect 30594 7736 30628 7770
rect 30594 7702 30628 7736
rect 30594 7668 30628 7702
rect 30594 7634 30628 7668
rect 30594 7600 30628 7634
rect 30594 7566 30628 7600
rect 30594 7532 30628 7566
rect 30594 7498 30628 7532
rect 30594 7464 30628 7498
rect 30594 7422 30628 7464
rect 30668 7422 30702 8398
rect 30796 7422 30830 8398
rect 30924 7422 30958 8398
rect 30998 8382 31032 8398
rect 30998 8348 31032 8382
rect 30998 8314 31032 8348
rect 30998 8280 31032 8314
rect 30998 8246 31032 8280
rect 30998 8212 31032 8246
rect 30998 8178 31032 8212
rect 30998 8144 31032 8178
rect 30998 8110 31032 8144
rect 30998 8076 31032 8110
rect 30998 8042 31032 8076
rect 30998 8008 31032 8042
rect 30998 7974 31032 8008
rect 30998 7940 31032 7974
rect 30998 7906 31032 7940
rect 30998 7872 31032 7906
rect 30998 7838 31032 7872
rect 30998 7804 31032 7838
rect 30998 7770 31032 7804
rect 30998 7736 31032 7770
rect 30998 7702 31032 7736
rect 30998 7668 31032 7702
rect 30998 7634 31032 7668
rect 30998 7600 31032 7634
rect 30998 7566 31032 7600
rect 30998 7532 31032 7566
rect 30998 7498 31032 7532
rect 30998 7464 31032 7498
rect 30998 7422 31032 7464
rect 31072 7422 31106 8398
rect 31200 7422 31234 8398
rect 31328 7422 31362 8398
rect 31402 8382 31436 8398
rect 31402 8348 31436 8382
rect 31402 8314 31436 8348
rect 31402 8280 31436 8314
rect 31402 8246 31436 8280
rect 31402 8212 31436 8246
rect 31402 8178 31436 8212
rect 31402 8144 31436 8178
rect 31402 8110 31436 8144
rect 31402 8076 31436 8110
rect 31402 8042 31436 8076
rect 31402 8008 31436 8042
rect 31402 7974 31436 8008
rect 31402 7940 31436 7974
rect 31402 7906 31436 7940
rect 31402 7872 31436 7906
rect 31402 7838 31436 7872
rect 31402 7804 31436 7838
rect 31402 7770 31436 7804
rect 31402 7736 31436 7770
rect 31402 7702 31436 7736
rect 31402 7668 31436 7702
rect 31402 7634 31436 7668
rect 31402 7600 31436 7634
rect 31402 7566 31436 7600
rect 31402 7532 31436 7566
rect 31402 7498 31436 7532
rect 31402 7464 31436 7498
rect 31402 7422 31436 7464
rect 746 7329 784 7363
rect 874 7329 912 7363
rect 1150 7329 1188 7363
rect 1278 7329 1316 7363
rect 1554 7329 1592 7363
rect 1682 7329 1720 7363
rect 1958 7329 1996 7363
rect 2086 7329 2124 7363
rect 2362 7329 2400 7363
rect 2490 7329 2528 7363
rect 2766 7329 2804 7363
rect 2894 7329 2932 7363
rect 7116 7329 7154 7363
rect 7244 7329 7282 7363
rect 7520 7329 7558 7363
rect 7648 7329 7686 7363
rect 7924 7329 7962 7363
rect 8052 7329 8090 7363
rect 8328 7329 8366 7363
rect 8456 7329 8494 7363
rect 8732 7329 8770 7363
rect 8860 7329 8898 7363
rect 9136 7329 9174 7363
rect 9264 7329 9302 7363
rect 13486 7329 13524 7363
rect 13614 7329 13652 7363
rect 13890 7329 13928 7363
rect 14018 7329 14056 7363
rect 14294 7329 14332 7363
rect 14422 7329 14460 7363
rect 14698 7329 14736 7363
rect 14826 7329 14864 7363
rect 15102 7329 15140 7363
rect 15230 7329 15268 7363
rect 15506 7329 15544 7363
rect 15634 7329 15672 7363
rect 19856 7329 19894 7363
rect 19984 7329 20022 7363
rect 20260 7329 20298 7363
rect 20388 7329 20426 7363
rect 20664 7329 20702 7363
rect 20792 7329 20830 7363
rect 21068 7329 21106 7363
rect 21196 7329 21234 7363
rect 21472 7329 21510 7363
rect 21600 7329 21638 7363
rect 21876 7329 21914 7363
rect 22004 7329 22042 7363
rect 29114 7329 29152 7363
rect 29242 7329 29280 7363
rect 29518 7329 29556 7363
rect 29646 7329 29684 7363
rect 29922 7329 29960 7363
rect 30050 7329 30088 7363
rect 30326 7329 30364 7363
rect 30454 7329 30492 7363
rect 30730 7329 30768 7363
rect 30858 7329 30896 7363
rect 31134 7329 31172 7363
rect 31262 7329 31300 7363
rect -4652 7279 -4614 7313
rect -4524 7279 -4486 7313
rect -4248 7279 -4210 7313
rect -4120 7279 -4082 7313
rect -3844 7279 -3806 7313
rect -3716 7279 -3678 7313
rect -3440 7279 -3402 7313
rect -3312 7279 -3274 7313
rect -3036 7279 -2998 7313
rect -2908 7279 -2870 7313
rect -2632 7279 -2594 7313
rect -2504 7279 -2466 7313
rect 935 6972 969 7006
rect 1029 6972 1063 7006
rect 1271 6972 1305 7006
rect 1365 6972 1399 7006
rect 1607 6972 1641 7006
rect 1701 6972 1735 7006
rect 1943 6972 1977 7006
rect 2037 6972 2071 7006
rect 2279 6972 2313 7006
rect 2373 6972 2407 7006
rect 2615 6972 2649 7006
rect 2709 6972 2743 7006
rect 7305 6972 7339 7006
rect 7399 6972 7433 7006
rect 7641 6972 7675 7006
rect 7735 6972 7769 7006
rect 7977 6972 8011 7006
rect 8071 6972 8105 7006
rect 8313 6972 8347 7006
rect 8407 6972 8441 7006
rect 8649 6972 8683 7006
rect 8743 6972 8777 7006
rect 8985 6972 9019 7006
rect 9079 6972 9113 7006
rect 13675 6972 13709 7006
rect 13769 6972 13803 7006
rect 14011 6972 14045 7006
rect 14105 6972 14139 7006
rect 14347 6972 14381 7006
rect 14441 6972 14475 7006
rect 14683 6972 14717 7006
rect 14777 6972 14811 7006
rect 15019 6972 15053 7006
rect 15113 6972 15147 7006
rect 15355 6972 15389 7006
rect 15449 6972 15483 7006
rect 20045 6972 20079 7006
rect 20139 6972 20173 7006
rect 20381 6972 20415 7006
rect 20475 6972 20509 7006
rect 20717 6972 20751 7006
rect 20811 6972 20845 7006
rect 21053 6972 21087 7006
rect 21147 6972 21181 7006
rect 21389 6972 21423 7006
rect 21483 6972 21517 7006
rect 21725 6972 21759 7006
rect 21819 6972 21853 7006
rect 29303 6972 29337 7006
rect 29397 6972 29431 7006
rect 29639 6972 29673 7006
rect 29733 6972 29767 7006
rect 29975 6972 30009 7006
rect 30069 6972 30103 7006
rect 30311 6972 30345 7006
rect 30405 6972 30439 7006
rect 30647 6972 30681 7006
rect 30741 6972 30775 7006
rect 30983 6972 31017 7006
rect 31077 6972 31111 7006
rect -4463 6922 -4429 6956
rect -4369 6922 -4335 6956
rect -4127 6922 -4093 6956
rect -4033 6922 -3999 6956
rect -3791 6922 -3757 6956
rect -3697 6922 -3663 6956
rect -3455 6922 -3421 6956
rect -3361 6922 -3327 6956
rect -3119 6922 -3085 6956
rect -3025 6922 -2991 6956
rect -2783 6922 -2749 6956
rect -2689 6922 -2655 6956
rect -4584 6830 -4550 6872
rect -4584 6796 -4550 6830
rect -4584 6762 -4550 6796
rect -4584 6728 -4550 6762
rect -4584 6694 -4550 6728
rect -4584 6660 -4550 6694
rect -4584 6626 -4550 6660
rect -4584 6592 -4550 6626
rect -4584 6558 -4550 6592
rect -4584 6524 -4550 6558
rect -4584 6490 -4550 6524
rect -4584 6456 -4550 6490
rect -4584 6422 -4550 6456
rect -4584 6388 -4550 6422
rect -4584 6354 -4550 6388
rect -4584 6320 -4550 6354
rect -4584 6286 -4550 6320
rect -4584 6252 -4550 6286
rect -4584 6218 -4550 6252
rect -4584 6184 -4550 6218
rect -4584 6150 -4550 6184
rect -4584 6116 -4550 6150
rect -4584 6082 -4550 6116
rect -4584 6048 -4550 6082
rect -4584 6014 -4550 6048
rect -4584 5980 -4550 6014
rect -4584 5946 -4550 5980
rect -4584 5912 -4550 5946
rect -4584 5896 -4550 5912
rect -4510 5896 -4476 6872
rect -4416 5896 -4382 6872
rect -4322 5896 -4288 6872
rect -4248 6856 -4214 6872
rect -4248 6822 -4214 6856
rect -4248 6788 -4214 6822
rect -4248 6754 -4214 6788
rect -4248 6720 -4214 6754
rect -4248 6686 -4214 6720
rect -4248 6652 -4214 6686
rect -4248 6618 -4214 6652
rect -4248 6584 -4214 6618
rect -4248 6550 -4214 6584
rect -4248 6516 -4214 6550
rect -4248 6482 -4214 6516
rect -4248 6448 -4214 6482
rect -4248 6414 -4214 6448
rect -4248 6380 -4214 6414
rect -4248 6346 -4214 6380
rect -4248 6312 -4214 6346
rect -4248 6278 -4214 6312
rect -4248 6244 -4214 6278
rect -4248 6210 -4214 6244
rect -4248 6176 -4214 6210
rect -4248 6142 -4214 6176
rect -4248 6108 -4214 6142
rect -4248 6074 -4214 6108
rect -4248 6040 -4214 6074
rect -4248 6006 -4214 6040
rect -4248 5972 -4214 6006
rect -4248 5938 -4214 5972
rect -4248 5896 -4214 5938
rect -4174 5896 -4140 6872
rect -4080 5896 -4046 6872
rect -3986 5896 -3952 6872
rect -3912 6856 -3878 6872
rect -3912 6822 -3878 6856
rect -3912 6788 -3878 6822
rect -3912 6754 -3878 6788
rect -3912 6720 -3878 6754
rect -3912 6686 -3878 6720
rect -3912 6652 -3878 6686
rect -3912 6618 -3878 6652
rect -3912 6584 -3878 6618
rect -3912 6550 -3878 6584
rect -3912 6516 -3878 6550
rect -3912 6482 -3878 6516
rect -3912 6448 -3878 6482
rect -3912 6414 -3878 6448
rect -3912 6380 -3878 6414
rect -3912 6346 -3878 6380
rect -3912 6312 -3878 6346
rect -3912 6278 -3878 6312
rect -3912 6244 -3878 6278
rect -3912 6210 -3878 6244
rect -3912 6176 -3878 6210
rect -3912 6142 -3878 6176
rect -3912 6108 -3878 6142
rect -3912 6074 -3878 6108
rect -3912 6040 -3878 6074
rect -3912 6006 -3878 6040
rect -3912 5972 -3878 6006
rect -3912 5938 -3878 5972
rect -3912 5896 -3878 5938
rect -3838 5896 -3804 6872
rect -3744 5896 -3710 6872
rect -3650 5896 -3616 6872
rect -3576 6856 -3542 6872
rect -3576 6822 -3542 6856
rect -3576 6788 -3542 6822
rect -3576 6754 -3542 6788
rect -3576 6720 -3542 6754
rect -3576 6686 -3542 6720
rect -3576 6652 -3542 6686
rect -3576 6618 -3542 6652
rect -3576 6584 -3542 6618
rect -3576 6550 -3542 6584
rect -3576 6516 -3542 6550
rect -3576 6482 -3542 6516
rect -3576 6448 -3542 6482
rect -3576 6414 -3542 6448
rect -3576 6380 -3542 6414
rect -3576 6346 -3542 6380
rect -3576 6312 -3542 6346
rect -3576 6278 -3542 6312
rect -3576 6244 -3542 6278
rect -3576 6210 -3542 6244
rect -3576 6176 -3542 6210
rect -3576 6142 -3542 6176
rect -3576 6108 -3542 6142
rect -3576 6074 -3542 6108
rect -3576 6040 -3542 6074
rect -3576 6006 -3542 6040
rect -3576 5972 -3542 6006
rect -3576 5938 -3542 5972
rect -3576 5896 -3542 5938
rect -3502 5896 -3468 6872
rect -3408 5896 -3374 6872
rect -3314 5896 -3280 6872
rect -3240 6856 -3206 6872
rect -3240 6822 -3206 6856
rect -3240 6788 -3206 6822
rect -3240 6754 -3206 6788
rect -3240 6720 -3206 6754
rect -3240 6686 -3206 6720
rect -3240 6652 -3206 6686
rect -3240 6618 -3206 6652
rect -3240 6584 -3206 6618
rect -3240 6550 -3206 6584
rect -3240 6516 -3206 6550
rect -3240 6482 -3206 6516
rect -3240 6448 -3206 6482
rect -3240 6414 -3206 6448
rect -3240 6380 -3206 6414
rect -3240 6346 -3206 6380
rect -3240 6312 -3206 6346
rect -3240 6278 -3206 6312
rect -3240 6244 -3206 6278
rect -3240 6210 -3206 6244
rect -3240 6176 -3206 6210
rect -3240 6142 -3206 6176
rect -3240 6108 -3206 6142
rect -3240 6074 -3206 6108
rect -3240 6040 -3206 6074
rect -3240 6006 -3206 6040
rect -3240 5972 -3206 6006
rect -3240 5938 -3206 5972
rect -3240 5896 -3206 5938
rect -3166 5896 -3132 6872
rect -3072 5896 -3038 6872
rect -2978 5896 -2944 6872
rect -2904 6856 -2870 6872
rect -2904 6822 -2870 6856
rect -2904 6788 -2870 6822
rect -2904 6754 -2870 6788
rect -2904 6720 -2870 6754
rect -2904 6686 -2870 6720
rect -2904 6652 -2870 6686
rect -2904 6618 -2870 6652
rect -2904 6584 -2870 6618
rect -2904 6550 -2870 6584
rect -2904 6516 -2870 6550
rect -2904 6482 -2870 6516
rect -2904 6448 -2870 6482
rect -2904 6414 -2870 6448
rect -2904 6380 -2870 6414
rect -2904 6346 -2870 6380
rect -2904 6312 -2870 6346
rect -2904 6278 -2870 6312
rect -2904 6244 -2870 6278
rect -2904 6210 -2870 6244
rect -2904 6176 -2870 6210
rect -2904 6142 -2870 6176
rect -2904 6108 -2870 6142
rect -2904 6074 -2870 6108
rect -2904 6040 -2870 6074
rect -2904 6006 -2870 6040
rect -2904 5972 -2870 6006
rect -2904 5938 -2870 5972
rect -2904 5896 -2870 5938
rect -2830 5896 -2796 6872
rect -2736 5896 -2702 6872
rect -2642 5896 -2608 6872
rect -2568 6856 -2534 6872
rect -2568 6822 -2534 6856
rect -2568 6788 -2534 6822
rect -2568 6754 -2534 6788
rect -2568 6720 -2534 6754
rect -2568 6686 -2534 6720
rect -2568 6652 -2534 6686
rect -2568 6618 -2534 6652
rect -2568 6584 -2534 6618
rect -2568 6550 -2534 6584
rect -2568 6516 -2534 6550
rect -2568 6482 -2534 6516
rect -2568 6448 -2534 6482
rect -2568 6414 -2534 6448
rect -2568 6380 -2534 6414
rect -2568 6346 -2534 6380
rect -2568 6312 -2534 6346
rect -2568 6278 -2534 6312
rect -2568 6244 -2534 6278
rect -2568 6210 -2534 6244
rect -2568 6176 -2534 6210
rect -2568 6142 -2534 6176
rect -2568 6108 -2534 6142
rect -2568 6074 -2534 6108
rect -2568 6040 -2534 6074
rect -2568 6006 -2534 6040
rect -2568 5972 -2534 6006
rect -2568 5938 -2534 5972
rect -2568 5896 -2534 5938
rect 814 6608 848 6634
rect 814 6574 848 6608
rect 814 6540 848 6574
rect 814 6506 848 6540
rect 814 6472 848 6506
rect 814 6438 848 6472
rect 814 6404 848 6438
rect 814 6370 848 6404
rect 814 6336 848 6370
rect 814 6302 848 6336
rect 814 6268 848 6302
rect 814 6234 848 6268
rect 814 6200 848 6234
rect 814 6166 848 6200
rect 814 6132 848 6166
rect 814 6098 848 6132
rect 814 6064 848 6098
rect 814 6030 848 6064
rect 814 5996 848 6030
rect 814 5962 848 5996
rect 814 5946 848 5962
rect 888 5946 922 6922
rect 982 5946 1016 6922
rect 1076 5946 1110 6922
rect 1150 6600 1184 6634
rect 1150 6566 1184 6600
rect 1150 6532 1184 6566
rect 1150 6498 1184 6532
rect 1150 6464 1184 6498
rect 1150 6430 1184 6464
rect 1150 6396 1184 6430
rect 1150 6362 1184 6396
rect 1150 6328 1184 6362
rect 1150 6294 1184 6328
rect 1150 6260 1184 6294
rect 1150 6226 1184 6260
rect 1150 6192 1184 6226
rect 1150 6158 1184 6192
rect 1150 6124 1184 6158
rect 1150 6090 1184 6124
rect 1150 6056 1184 6090
rect 1150 6022 1184 6056
rect 1150 5988 1184 6022
rect 1150 5946 1184 5988
rect 1224 5946 1258 6922
rect 1318 5946 1352 6922
rect 1412 5946 1446 6922
rect 1486 6600 1520 6634
rect 1486 6566 1520 6600
rect 1486 6532 1520 6566
rect 1486 6498 1520 6532
rect 1486 6464 1520 6498
rect 1486 6430 1520 6464
rect 1486 6396 1520 6430
rect 1486 6362 1520 6396
rect 1486 6328 1520 6362
rect 1486 6294 1520 6328
rect 1486 6260 1520 6294
rect 1486 6226 1520 6260
rect 1486 6192 1520 6226
rect 1486 6158 1520 6192
rect 1486 6124 1520 6158
rect 1486 6090 1520 6124
rect 1486 6056 1520 6090
rect 1486 6022 1520 6056
rect 1486 5988 1520 6022
rect 1486 5946 1520 5988
rect 1560 5946 1594 6922
rect 1654 5946 1688 6922
rect 1748 5946 1782 6922
rect 1822 6600 1856 6634
rect 1822 6566 1856 6600
rect 1822 6532 1856 6566
rect 1822 6498 1856 6532
rect 1822 6464 1856 6498
rect 1822 6430 1856 6464
rect 1822 6396 1856 6430
rect 1822 6362 1856 6396
rect 1822 6328 1856 6362
rect 1822 6294 1856 6328
rect 1822 6260 1856 6294
rect 1822 6226 1856 6260
rect 1822 6192 1856 6226
rect 1822 6158 1856 6192
rect 1822 6124 1856 6158
rect 1822 6090 1856 6124
rect 1822 6056 1856 6090
rect 1822 6022 1856 6056
rect 1822 5988 1856 6022
rect 1822 5946 1856 5988
rect 1896 5946 1930 6922
rect 1990 5946 2024 6922
rect 2084 5946 2118 6922
rect 2158 6600 2192 6634
rect 2158 6566 2192 6600
rect 2158 6532 2192 6566
rect 2158 6498 2192 6532
rect 2158 6464 2192 6498
rect 2158 6430 2192 6464
rect 2158 6396 2192 6430
rect 2158 6362 2192 6396
rect 2158 6328 2192 6362
rect 2158 6294 2192 6328
rect 2158 6260 2192 6294
rect 2158 6226 2192 6260
rect 2158 6192 2192 6226
rect 2158 6158 2192 6192
rect 2158 6124 2192 6158
rect 2158 6090 2192 6124
rect 2158 6056 2192 6090
rect 2158 6022 2192 6056
rect 2158 5988 2192 6022
rect 2158 5946 2192 5988
rect 2232 5946 2266 6922
rect 2326 5946 2360 6922
rect 2420 5946 2454 6922
rect 2494 6600 2528 6634
rect 2494 6566 2528 6600
rect 2494 6532 2528 6566
rect 2494 6498 2528 6532
rect 2494 6464 2528 6498
rect 2494 6430 2528 6464
rect 2494 6396 2528 6430
rect 2494 6362 2528 6396
rect 2494 6328 2528 6362
rect 2494 6294 2528 6328
rect 2494 6260 2528 6294
rect 2494 6226 2528 6260
rect 2494 6192 2528 6226
rect 2494 6158 2528 6192
rect 2494 6124 2528 6158
rect 2494 6090 2528 6124
rect 2494 6056 2528 6090
rect 2494 6022 2528 6056
rect 2494 5988 2528 6022
rect 2494 5946 2528 5988
rect 2568 5946 2602 6922
rect 2662 5946 2696 6922
rect 2756 5946 2790 6922
rect 2830 6600 2864 6634
rect 2830 6566 2864 6600
rect 2830 6532 2864 6566
rect 2830 6498 2864 6532
rect 2830 6464 2864 6498
rect 2830 6430 2864 6464
rect 2830 6396 2864 6430
rect 2830 6362 2864 6396
rect 2830 6328 2864 6362
rect 2830 6294 2864 6328
rect 2830 6260 2864 6294
rect 2830 6226 2864 6260
rect 2830 6192 2864 6226
rect 2830 6158 2864 6192
rect 2830 6124 2864 6158
rect 2830 6090 2864 6124
rect 2830 6056 2864 6090
rect 2830 6022 2864 6056
rect 2830 5988 2864 6022
rect 2830 5946 2864 5988
rect 7184 6608 7218 6634
rect 7184 6574 7218 6608
rect 7184 6540 7218 6574
rect 7184 6506 7218 6540
rect 7184 6472 7218 6506
rect 7184 6438 7218 6472
rect 7184 6404 7218 6438
rect 7184 6370 7218 6404
rect 7184 6336 7218 6370
rect 7184 6302 7218 6336
rect 7184 6268 7218 6302
rect 7184 6234 7218 6268
rect 7184 6200 7218 6234
rect 7184 6166 7218 6200
rect 7184 6132 7218 6166
rect 7184 6098 7218 6132
rect 7184 6064 7218 6098
rect 7184 6030 7218 6064
rect 7184 5996 7218 6030
rect 7184 5962 7218 5996
rect 7184 5946 7218 5962
rect 7258 5946 7292 6922
rect 7352 5946 7386 6922
rect 7446 5946 7480 6922
rect 7520 6600 7554 6634
rect 7520 6566 7554 6600
rect 7520 6532 7554 6566
rect 7520 6498 7554 6532
rect 7520 6464 7554 6498
rect 7520 6430 7554 6464
rect 7520 6396 7554 6430
rect 7520 6362 7554 6396
rect 7520 6328 7554 6362
rect 7520 6294 7554 6328
rect 7520 6260 7554 6294
rect 7520 6226 7554 6260
rect 7520 6192 7554 6226
rect 7520 6158 7554 6192
rect 7520 6124 7554 6158
rect 7520 6090 7554 6124
rect 7520 6056 7554 6090
rect 7520 6022 7554 6056
rect 7520 5988 7554 6022
rect 7520 5946 7554 5988
rect 7594 5946 7628 6922
rect 7688 5946 7722 6922
rect 7782 5946 7816 6922
rect 7856 6600 7890 6634
rect 7856 6566 7890 6600
rect 7856 6532 7890 6566
rect 7856 6498 7890 6532
rect 7856 6464 7890 6498
rect 7856 6430 7890 6464
rect 7856 6396 7890 6430
rect 7856 6362 7890 6396
rect 7856 6328 7890 6362
rect 7856 6294 7890 6328
rect 7856 6260 7890 6294
rect 7856 6226 7890 6260
rect 7856 6192 7890 6226
rect 7856 6158 7890 6192
rect 7856 6124 7890 6158
rect 7856 6090 7890 6124
rect 7856 6056 7890 6090
rect 7856 6022 7890 6056
rect 7856 5988 7890 6022
rect 7856 5946 7890 5988
rect 7930 5946 7964 6922
rect 8024 5946 8058 6922
rect 8118 5946 8152 6922
rect 8192 6600 8226 6634
rect 8192 6566 8226 6600
rect 8192 6532 8226 6566
rect 8192 6498 8226 6532
rect 8192 6464 8226 6498
rect 8192 6430 8226 6464
rect 8192 6396 8226 6430
rect 8192 6362 8226 6396
rect 8192 6328 8226 6362
rect 8192 6294 8226 6328
rect 8192 6260 8226 6294
rect 8192 6226 8226 6260
rect 8192 6192 8226 6226
rect 8192 6158 8226 6192
rect 8192 6124 8226 6158
rect 8192 6090 8226 6124
rect 8192 6056 8226 6090
rect 8192 6022 8226 6056
rect 8192 5988 8226 6022
rect 8192 5946 8226 5988
rect 8266 5946 8300 6922
rect 8360 5946 8394 6922
rect 8454 5946 8488 6922
rect 8528 6600 8562 6634
rect 8528 6566 8562 6600
rect 8528 6532 8562 6566
rect 8528 6498 8562 6532
rect 8528 6464 8562 6498
rect 8528 6430 8562 6464
rect 8528 6396 8562 6430
rect 8528 6362 8562 6396
rect 8528 6328 8562 6362
rect 8528 6294 8562 6328
rect 8528 6260 8562 6294
rect 8528 6226 8562 6260
rect 8528 6192 8562 6226
rect 8528 6158 8562 6192
rect 8528 6124 8562 6158
rect 8528 6090 8562 6124
rect 8528 6056 8562 6090
rect 8528 6022 8562 6056
rect 8528 5988 8562 6022
rect 8528 5946 8562 5988
rect 8602 5946 8636 6922
rect 8696 5946 8730 6922
rect 8790 5946 8824 6922
rect 8864 6600 8898 6634
rect 8864 6566 8898 6600
rect 8864 6532 8898 6566
rect 8864 6498 8898 6532
rect 8864 6464 8898 6498
rect 8864 6430 8898 6464
rect 8864 6396 8898 6430
rect 8864 6362 8898 6396
rect 8864 6328 8898 6362
rect 8864 6294 8898 6328
rect 8864 6260 8898 6294
rect 8864 6226 8898 6260
rect 8864 6192 8898 6226
rect 8864 6158 8898 6192
rect 8864 6124 8898 6158
rect 8864 6090 8898 6124
rect 8864 6056 8898 6090
rect 8864 6022 8898 6056
rect 8864 5988 8898 6022
rect 8864 5946 8898 5988
rect 8938 5946 8972 6922
rect 9032 5946 9066 6922
rect 9126 5946 9160 6922
rect 9200 6600 9234 6634
rect 9200 6566 9234 6600
rect 9200 6532 9234 6566
rect 9200 6498 9234 6532
rect 9200 6464 9234 6498
rect 9200 6430 9234 6464
rect 9200 6396 9234 6430
rect 9200 6362 9234 6396
rect 9200 6328 9234 6362
rect 9200 6294 9234 6328
rect 9200 6260 9234 6294
rect 9200 6226 9234 6260
rect 9200 6192 9234 6226
rect 9200 6158 9234 6192
rect 9200 6124 9234 6158
rect 9200 6090 9234 6124
rect 9200 6056 9234 6090
rect 9200 6022 9234 6056
rect 9200 5988 9234 6022
rect 9200 5946 9234 5988
rect 13554 6608 13588 6634
rect 13554 6574 13588 6608
rect 13554 6540 13588 6574
rect 13554 6506 13588 6540
rect 13554 6472 13588 6506
rect 13554 6438 13588 6472
rect 13554 6404 13588 6438
rect 13554 6370 13588 6404
rect 13554 6336 13588 6370
rect 13554 6302 13588 6336
rect 13554 6268 13588 6302
rect 13554 6234 13588 6268
rect 13554 6200 13588 6234
rect 13554 6166 13588 6200
rect 13554 6132 13588 6166
rect 13554 6098 13588 6132
rect 13554 6064 13588 6098
rect 13554 6030 13588 6064
rect 13554 5996 13588 6030
rect 13554 5962 13588 5996
rect 13554 5946 13588 5962
rect 13628 5946 13662 6922
rect 13722 5946 13756 6922
rect 13816 5946 13850 6922
rect 13890 6600 13924 6634
rect 13890 6566 13924 6600
rect 13890 6532 13924 6566
rect 13890 6498 13924 6532
rect 13890 6464 13924 6498
rect 13890 6430 13924 6464
rect 13890 6396 13924 6430
rect 13890 6362 13924 6396
rect 13890 6328 13924 6362
rect 13890 6294 13924 6328
rect 13890 6260 13924 6294
rect 13890 6226 13924 6260
rect 13890 6192 13924 6226
rect 13890 6158 13924 6192
rect 13890 6124 13924 6158
rect 13890 6090 13924 6124
rect 13890 6056 13924 6090
rect 13890 6022 13924 6056
rect 13890 5988 13924 6022
rect 13890 5946 13924 5988
rect 13964 5946 13998 6922
rect 14058 5946 14092 6922
rect 14152 5946 14186 6922
rect 14226 6600 14260 6634
rect 14226 6566 14260 6600
rect 14226 6532 14260 6566
rect 14226 6498 14260 6532
rect 14226 6464 14260 6498
rect 14226 6430 14260 6464
rect 14226 6396 14260 6430
rect 14226 6362 14260 6396
rect 14226 6328 14260 6362
rect 14226 6294 14260 6328
rect 14226 6260 14260 6294
rect 14226 6226 14260 6260
rect 14226 6192 14260 6226
rect 14226 6158 14260 6192
rect 14226 6124 14260 6158
rect 14226 6090 14260 6124
rect 14226 6056 14260 6090
rect 14226 6022 14260 6056
rect 14226 5988 14260 6022
rect 14226 5946 14260 5988
rect 14300 5946 14334 6922
rect 14394 5946 14428 6922
rect 14488 5946 14522 6922
rect 14562 6600 14596 6634
rect 14562 6566 14596 6600
rect 14562 6532 14596 6566
rect 14562 6498 14596 6532
rect 14562 6464 14596 6498
rect 14562 6430 14596 6464
rect 14562 6396 14596 6430
rect 14562 6362 14596 6396
rect 14562 6328 14596 6362
rect 14562 6294 14596 6328
rect 14562 6260 14596 6294
rect 14562 6226 14596 6260
rect 14562 6192 14596 6226
rect 14562 6158 14596 6192
rect 14562 6124 14596 6158
rect 14562 6090 14596 6124
rect 14562 6056 14596 6090
rect 14562 6022 14596 6056
rect 14562 5988 14596 6022
rect 14562 5946 14596 5988
rect 14636 5946 14670 6922
rect 14730 5946 14764 6922
rect 14824 5946 14858 6922
rect 14898 6600 14932 6634
rect 14898 6566 14932 6600
rect 14898 6532 14932 6566
rect 14898 6498 14932 6532
rect 14898 6464 14932 6498
rect 14898 6430 14932 6464
rect 14898 6396 14932 6430
rect 14898 6362 14932 6396
rect 14898 6328 14932 6362
rect 14898 6294 14932 6328
rect 14898 6260 14932 6294
rect 14898 6226 14932 6260
rect 14898 6192 14932 6226
rect 14898 6158 14932 6192
rect 14898 6124 14932 6158
rect 14898 6090 14932 6124
rect 14898 6056 14932 6090
rect 14898 6022 14932 6056
rect 14898 5988 14932 6022
rect 14898 5946 14932 5988
rect 14972 5946 15006 6922
rect 15066 5946 15100 6922
rect 15160 5946 15194 6922
rect 15234 6600 15268 6634
rect 15234 6566 15268 6600
rect 15234 6532 15268 6566
rect 15234 6498 15268 6532
rect 15234 6464 15268 6498
rect 15234 6430 15268 6464
rect 15234 6396 15268 6430
rect 15234 6362 15268 6396
rect 15234 6328 15268 6362
rect 15234 6294 15268 6328
rect 15234 6260 15268 6294
rect 15234 6226 15268 6260
rect 15234 6192 15268 6226
rect 15234 6158 15268 6192
rect 15234 6124 15268 6158
rect 15234 6090 15268 6124
rect 15234 6056 15268 6090
rect 15234 6022 15268 6056
rect 15234 5988 15268 6022
rect 15234 5946 15268 5988
rect 15308 5946 15342 6922
rect 15402 5946 15436 6922
rect 15496 5946 15530 6922
rect 15570 6600 15604 6634
rect 15570 6566 15604 6600
rect 15570 6532 15604 6566
rect 15570 6498 15604 6532
rect 15570 6464 15604 6498
rect 15570 6430 15604 6464
rect 15570 6396 15604 6430
rect 15570 6362 15604 6396
rect 15570 6328 15604 6362
rect 15570 6294 15604 6328
rect 15570 6260 15604 6294
rect 15570 6226 15604 6260
rect 15570 6192 15604 6226
rect 15570 6158 15604 6192
rect 15570 6124 15604 6158
rect 15570 6090 15604 6124
rect 15570 6056 15604 6090
rect 15570 6022 15604 6056
rect 15570 5988 15604 6022
rect 15570 5946 15604 5988
rect 19924 6608 19958 6634
rect 19924 6574 19958 6608
rect 19924 6540 19958 6574
rect 19924 6506 19958 6540
rect 19924 6472 19958 6506
rect 19924 6438 19958 6472
rect 19924 6404 19958 6438
rect 19924 6370 19958 6404
rect 19924 6336 19958 6370
rect 19924 6302 19958 6336
rect 19924 6268 19958 6302
rect 19924 6234 19958 6268
rect 19924 6200 19958 6234
rect 19924 6166 19958 6200
rect 19924 6132 19958 6166
rect 19924 6098 19958 6132
rect 19924 6064 19958 6098
rect 19924 6030 19958 6064
rect 19924 5996 19958 6030
rect 19924 5962 19958 5996
rect 19924 5946 19958 5962
rect 19998 5946 20032 6922
rect 20092 5946 20126 6922
rect 20186 5946 20220 6922
rect 20260 6600 20294 6634
rect 20260 6566 20294 6600
rect 20260 6532 20294 6566
rect 20260 6498 20294 6532
rect 20260 6464 20294 6498
rect 20260 6430 20294 6464
rect 20260 6396 20294 6430
rect 20260 6362 20294 6396
rect 20260 6328 20294 6362
rect 20260 6294 20294 6328
rect 20260 6260 20294 6294
rect 20260 6226 20294 6260
rect 20260 6192 20294 6226
rect 20260 6158 20294 6192
rect 20260 6124 20294 6158
rect 20260 6090 20294 6124
rect 20260 6056 20294 6090
rect 20260 6022 20294 6056
rect 20260 5988 20294 6022
rect 20260 5946 20294 5988
rect 20334 5946 20368 6922
rect 20428 5946 20462 6922
rect 20522 5946 20556 6922
rect 20596 6600 20630 6634
rect 20596 6566 20630 6600
rect 20596 6532 20630 6566
rect 20596 6498 20630 6532
rect 20596 6464 20630 6498
rect 20596 6430 20630 6464
rect 20596 6396 20630 6430
rect 20596 6362 20630 6396
rect 20596 6328 20630 6362
rect 20596 6294 20630 6328
rect 20596 6260 20630 6294
rect 20596 6226 20630 6260
rect 20596 6192 20630 6226
rect 20596 6158 20630 6192
rect 20596 6124 20630 6158
rect 20596 6090 20630 6124
rect 20596 6056 20630 6090
rect 20596 6022 20630 6056
rect 20596 5988 20630 6022
rect 20596 5946 20630 5988
rect 20670 5946 20704 6922
rect 20764 5946 20798 6922
rect 20858 5946 20892 6922
rect 20932 6600 20966 6634
rect 20932 6566 20966 6600
rect 20932 6532 20966 6566
rect 20932 6498 20966 6532
rect 20932 6464 20966 6498
rect 20932 6430 20966 6464
rect 20932 6396 20966 6430
rect 20932 6362 20966 6396
rect 20932 6328 20966 6362
rect 20932 6294 20966 6328
rect 20932 6260 20966 6294
rect 20932 6226 20966 6260
rect 20932 6192 20966 6226
rect 20932 6158 20966 6192
rect 20932 6124 20966 6158
rect 20932 6090 20966 6124
rect 20932 6056 20966 6090
rect 20932 6022 20966 6056
rect 20932 5988 20966 6022
rect 20932 5946 20966 5988
rect 21006 5946 21040 6922
rect 21100 5946 21134 6922
rect 21194 5946 21228 6922
rect 21268 6600 21302 6634
rect 21268 6566 21302 6600
rect 21268 6532 21302 6566
rect 21268 6498 21302 6532
rect 21268 6464 21302 6498
rect 21268 6430 21302 6464
rect 21268 6396 21302 6430
rect 21268 6362 21302 6396
rect 21268 6328 21302 6362
rect 21268 6294 21302 6328
rect 21268 6260 21302 6294
rect 21268 6226 21302 6260
rect 21268 6192 21302 6226
rect 21268 6158 21302 6192
rect 21268 6124 21302 6158
rect 21268 6090 21302 6124
rect 21268 6056 21302 6090
rect 21268 6022 21302 6056
rect 21268 5988 21302 6022
rect 21268 5946 21302 5988
rect 21342 5946 21376 6922
rect 21436 5946 21470 6922
rect 21530 5946 21564 6922
rect 21604 6600 21638 6634
rect 21604 6566 21638 6600
rect 21604 6532 21638 6566
rect 21604 6498 21638 6532
rect 21604 6464 21638 6498
rect 21604 6430 21638 6464
rect 21604 6396 21638 6430
rect 21604 6362 21638 6396
rect 21604 6328 21638 6362
rect 21604 6294 21638 6328
rect 21604 6260 21638 6294
rect 21604 6226 21638 6260
rect 21604 6192 21638 6226
rect 21604 6158 21638 6192
rect 21604 6124 21638 6158
rect 21604 6090 21638 6124
rect 21604 6056 21638 6090
rect 21604 6022 21638 6056
rect 21604 5988 21638 6022
rect 21604 5946 21638 5988
rect 21678 5946 21712 6922
rect 21772 5946 21806 6922
rect 21866 5946 21900 6922
rect 21940 6600 21974 6634
rect 21940 6566 21974 6600
rect 21940 6532 21974 6566
rect 21940 6498 21974 6532
rect 21940 6464 21974 6498
rect 21940 6430 21974 6464
rect 21940 6396 21974 6430
rect 21940 6362 21974 6396
rect 21940 6328 21974 6362
rect 21940 6294 21974 6328
rect 21940 6260 21974 6294
rect 21940 6226 21974 6260
rect 21940 6192 21974 6226
rect 21940 6158 21974 6192
rect 21940 6124 21974 6158
rect 21940 6090 21974 6124
rect 21940 6056 21974 6090
rect 21940 6022 21974 6056
rect 21940 5988 21974 6022
rect 21940 5946 21974 5988
rect 29182 6608 29216 6634
rect 29182 6574 29216 6608
rect 29182 6540 29216 6574
rect 29182 6506 29216 6540
rect 29182 6472 29216 6506
rect 29182 6438 29216 6472
rect 29182 6404 29216 6438
rect 29182 6370 29216 6404
rect 29182 6336 29216 6370
rect 29182 6302 29216 6336
rect 29182 6268 29216 6302
rect 29182 6234 29216 6268
rect 29182 6200 29216 6234
rect 29182 6166 29216 6200
rect 29182 6132 29216 6166
rect 29182 6098 29216 6132
rect 29182 6064 29216 6098
rect 29182 6030 29216 6064
rect 29182 5996 29216 6030
rect 29182 5962 29216 5996
rect 29182 5946 29216 5962
rect 29256 5946 29290 6922
rect 29350 5946 29384 6922
rect 29444 5946 29478 6922
rect 29518 6600 29552 6634
rect 29518 6566 29552 6600
rect 29518 6532 29552 6566
rect 29518 6498 29552 6532
rect 29518 6464 29552 6498
rect 29518 6430 29552 6464
rect 29518 6396 29552 6430
rect 29518 6362 29552 6396
rect 29518 6328 29552 6362
rect 29518 6294 29552 6328
rect 29518 6260 29552 6294
rect 29518 6226 29552 6260
rect 29518 6192 29552 6226
rect 29518 6158 29552 6192
rect 29518 6124 29552 6158
rect 29518 6090 29552 6124
rect 29518 6056 29552 6090
rect 29518 6022 29552 6056
rect 29518 5988 29552 6022
rect 29518 5946 29552 5988
rect 29592 5946 29626 6922
rect 29686 5946 29720 6922
rect 29780 5946 29814 6922
rect 29854 6600 29888 6634
rect 29854 6566 29888 6600
rect 29854 6532 29888 6566
rect 29854 6498 29888 6532
rect 29854 6464 29888 6498
rect 29854 6430 29888 6464
rect 29854 6396 29888 6430
rect 29854 6362 29888 6396
rect 29854 6328 29888 6362
rect 29854 6294 29888 6328
rect 29854 6260 29888 6294
rect 29854 6226 29888 6260
rect 29854 6192 29888 6226
rect 29854 6158 29888 6192
rect 29854 6124 29888 6158
rect 29854 6090 29888 6124
rect 29854 6056 29888 6090
rect 29854 6022 29888 6056
rect 29854 5988 29888 6022
rect 29854 5946 29888 5988
rect 29928 5946 29962 6922
rect 30022 5946 30056 6922
rect 30116 5946 30150 6922
rect 30190 6600 30224 6634
rect 30190 6566 30224 6600
rect 30190 6532 30224 6566
rect 30190 6498 30224 6532
rect 30190 6464 30224 6498
rect 30190 6430 30224 6464
rect 30190 6396 30224 6430
rect 30190 6362 30224 6396
rect 30190 6328 30224 6362
rect 30190 6294 30224 6328
rect 30190 6260 30224 6294
rect 30190 6226 30224 6260
rect 30190 6192 30224 6226
rect 30190 6158 30224 6192
rect 30190 6124 30224 6158
rect 30190 6090 30224 6124
rect 30190 6056 30224 6090
rect 30190 6022 30224 6056
rect 30190 5988 30224 6022
rect 30190 5946 30224 5988
rect 30264 5946 30298 6922
rect 30358 5946 30392 6922
rect 30452 5946 30486 6922
rect 30526 6600 30560 6634
rect 30526 6566 30560 6600
rect 30526 6532 30560 6566
rect 30526 6498 30560 6532
rect 30526 6464 30560 6498
rect 30526 6430 30560 6464
rect 30526 6396 30560 6430
rect 30526 6362 30560 6396
rect 30526 6328 30560 6362
rect 30526 6294 30560 6328
rect 30526 6260 30560 6294
rect 30526 6226 30560 6260
rect 30526 6192 30560 6226
rect 30526 6158 30560 6192
rect 30526 6124 30560 6158
rect 30526 6090 30560 6124
rect 30526 6056 30560 6090
rect 30526 6022 30560 6056
rect 30526 5988 30560 6022
rect 30526 5946 30560 5988
rect 30600 5946 30634 6922
rect 30694 5946 30728 6922
rect 30788 5946 30822 6922
rect 30862 6600 30896 6634
rect 30862 6566 30896 6600
rect 30862 6532 30896 6566
rect 30862 6498 30896 6532
rect 30862 6464 30896 6498
rect 30862 6430 30896 6464
rect 30862 6396 30896 6430
rect 30862 6362 30896 6396
rect 30862 6328 30896 6362
rect 30862 6294 30896 6328
rect 30862 6260 30896 6294
rect 30862 6226 30896 6260
rect 30862 6192 30896 6226
rect 30862 6158 30896 6192
rect 30862 6124 30896 6158
rect 30862 6090 30896 6124
rect 30862 6056 30896 6090
rect 30862 6022 30896 6056
rect 30862 5988 30896 6022
rect 30862 5946 30896 5988
rect 30936 5946 30970 6922
rect 31030 5946 31064 6922
rect 31124 5946 31158 6922
rect 31198 6600 31232 6634
rect 31198 6566 31232 6600
rect 31198 6532 31232 6566
rect 31198 6498 31232 6532
rect 31198 6464 31232 6498
rect 31198 6430 31232 6464
rect 31198 6396 31232 6430
rect 31198 6362 31232 6396
rect 31198 6328 31232 6362
rect 31198 6294 31232 6328
rect 31198 6260 31232 6294
rect 31198 6226 31232 6260
rect 31198 6192 31232 6226
rect 31198 6158 31232 6192
rect 31198 6124 31232 6158
rect 31198 6090 31232 6124
rect 31198 6056 31232 6090
rect 31198 6022 31232 6056
rect 31198 5988 31232 6022
rect 31198 5946 31232 5988
rect -4463 5812 -4429 5846
rect -4369 5812 -4335 5846
rect -4127 5812 -4093 5846
rect -4033 5812 -3999 5846
rect -3791 5812 -3757 5846
rect -3697 5812 -3663 5846
rect -3455 5812 -3421 5846
rect -3361 5812 -3327 5846
rect -3119 5812 -3085 5846
rect -3025 5812 -2991 5846
rect -2783 5812 -2749 5846
rect -2689 5812 -2655 5846
<< metal1 >>
rect 450 8872 562 8882
rect -4948 8822 -4836 8832
rect -4948 8654 -4918 8822
rect -4862 8654 -4836 8822
rect -5242 6616 -4984 8522
rect -4948 7072 -4836 8654
rect 450 8704 480 8872
rect 536 8704 562 8872
rect -4808 8552 -2312 8558
rect -4808 8500 -4788 8552
rect -4808 8494 -2312 8500
rect -4808 8360 -4696 8494
rect -4666 8441 -4472 8448
rect -4666 8407 -4652 8441
rect -4614 8407 -4524 8441
rect -4486 8407 -4472 8441
rect -4666 8400 -4472 8407
rect -4424 8360 -4312 8494
rect -4262 8441 -4068 8448
rect -4262 8407 -4248 8441
rect -4210 8407 -4120 8441
rect -4082 8407 -4068 8441
rect -4262 8400 -4068 8407
rect -4020 8360 -3908 8494
rect -3858 8441 -3664 8448
rect -3858 8407 -3844 8441
rect -3806 8407 -3716 8441
rect -3678 8407 -3664 8441
rect -3858 8400 -3664 8407
rect -3616 8360 -3504 8494
rect -3454 8441 -3260 8448
rect -3454 8407 -3440 8441
rect -3402 8407 -3312 8441
rect -3274 8407 -3260 8441
rect -3454 8400 -3260 8407
rect -3212 8360 -3100 8494
rect -3050 8441 -2856 8448
rect -3050 8407 -3036 8441
rect -2998 8407 -2908 8441
rect -2870 8407 -2856 8441
rect -3050 8400 -2856 8407
rect -2808 8360 -2696 8494
rect -2646 8441 -2452 8448
rect -2646 8407 -2632 8441
rect -2594 8407 -2504 8441
rect -2466 8407 -2452 8441
rect -2646 8400 -2452 8407
rect -2424 8360 -2312 8494
rect -4808 8348 -4674 8360
rect -4592 8358 -4546 8360
rect -4808 7372 -4788 8348
rect -4754 7372 -4714 8348
rect -4680 7372 -4674 8348
rect -4808 7360 -4674 7372
rect -4598 8348 -4540 8358
rect -4598 7366 -4540 7372
rect -4464 8348 -4270 8360
rect -4188 8358 -4142 8360
rect -4464 7372 -4458 8348
rect -4424 7372 -4384 8348
rect -4350 7372 -4310 8348
rect -4276 7372 -4270 8348
rect -4592 7360 -4546 7366
rect -4464 7360 -4270 7372
rect -4194 8348 -4136 8358
rect -4194 7366 -4136 7372
rect -4060 8348 -3866 8360
rect -3784 8358 -3738 8360
rect -4060 7372 -4054 8348
rect -4020 7372 -3980 8348
rect -3946 7372 -3906 8348
rect -3872 7372 -3866 8348
rect -4188 7360 -4142 7366
rect -4060 7360 -3866 7372
rect -3790 8348 -3732 8358
rect -3790 7366 -3732 7372
rect -3656 8348 -3462 8360
rect -3380 8358 -3334 8360
rect -3656 7372 -3650 8348
rect -3616 7372 -3576 8348
rect -3542 7372 -3502 8348
rect -3468 7372 -3462 8348
rect -3784 7360 -3738 7366
rect -3656 7360 -3462 7372
rect -3386 8348 -3328 8358
rect -3386 7366 -3328 7372
rect -3252 8348 -3058 8360
rect -2976 8358 -2930 8360
rect -3252 7372 -3246 8348
rect -3212 7372 -3172 8348
rect -3138 7372 -3098 8348
rect -3064 7372 -3058 8348
rect -3380 7360 -3334 7366
rect -3252 7360 -3058 7372
rect -2982 8348 -2924 8358
rect -2982 7366 -2924 7372
rect -2848 8348 -2654 8360
rect -2572 8358 -2526 8360
rect -2848 7372 -2842 8348
rect -2808 7372 -2768 8348
rect -2734 7372 -2694 8348
rect -2660 7372 -2654 8348
rect -2976 7360 -2930 7366
rect -2848 7360 -2654 7372
rect -2578 8348 -2520 8358
rect -2578 7366 -2520 7372
rect -2444 8348 -2312 8360
rect -2444 7372 -2438 8348
rect -2404 7372 -2364 8348
rect -2330 7372 -2312 8348
rect -2572 7360 -2526 7366
rect -2444 7360 -2312 7372
rect -4666 7313 -4472 7320
rect -4666 7279 -4652 7313
rect -4614 7279 -4524 7313
rect -4486 7279 -4472 7313
rect -4666 7260 -4472 7279
rect -4262 7313 -4068 7320
rect -4262 7279 -4248 7313
rect -4210 7279 -4120 7313
rect -4082 7279 -4068 7313
rect -4262 7260 -4068 7279
rect -3858 7313 -3664 7320
rect -3858 7279 -3844 7313
rect -3806 7279 -3716 7313
rect -3678 7279 -3664 7313
rect -4594 7218 -4472 7260
rect -4594 7212 -4344 7218
rect -4370 7160 -4344 7212
rect -4594 7154 -4344 7160
rect -4948 7014 -4836 7020
rect -4478 6972 -4344 7154
rect -4232 7078 -4098 7260
rect -3858 7218 -3664 7279
rect -3454 7313 -3260 7320
rect -3454 7279 -3440 7313
rect -3402 7279 -3312 7313
rect -3274 7279 -3260 7313
rect -3858 7212 -3634 7218
rect -3858 7154 -3634 7160
rect -4232 7072 -3984 7078
rect -4008 7020 -3984 7072
rect -4232 7014 -3984 7020
rect -4478 6956 -4320 6972
rect -4478 6922 -4463 6956
rect -4429 6922 -4369 6956
rect -4335 6922 -4320 6956
rect -4478 6916 -4320 6922
rect -4142 6956 -3984 7014
rect -4142 6922 -4127 6956
rect -4093 6922 -4033 6956
rect -3999 6922 -3984 6956
rect -4142 6916 -3984 6922
rect -3806 6956 -3648 7154
rect -3454 7078 -3260 7279
rect -3050 7313 -2856 7320
rect -3050 7279 -3036 7313
rect -2998 7279 -2908 7313
rect -2870 7279 -2856 7313
rect -3050 7218 -2856 7279
rect -3104 7212 -2856 7218
rect -2880 7160 -2856 7212
rect -3104 7154 -2856 7160
rect -2646 7313 -2452 7320
rect -2646 7279 -2632 7313
rect -2594 7279 -2504 7313
rect -2466 7279 -2452 7313
rect -2646 7242 -2452 7279
rect -3478 7072 -3254 7078
rect -3478 7014 -3254 7020
rect -3806 6922 -3791 6956
rect -3757 6922 -3697 6956
rect -3663 6922 -3648 6956
rect -3806 6916 -3648 6922
rect -3470 6956 -3312 7014
rect -3104 6972 -2992 7154
rect -2646 7078 -2526 7242
rect -2758 7072 -2526 7078
rect -2534 7020 -2526 7072
rect -2758 7014 -2526 7020
rect -2418 7212 -2306 7218
rect -2758 6972 -2640 7014
rect -3470 6922 -3455 6956
rect -3421 6922 -3361 6956
rect -3327 6922 -3312 6956
rect -3470 6916 -3312 6922
rect -3134 6956 -2976 6972
rect -3134 6922 -3119 6956
rect -3085 6922 -3025 6956
rect -2991 6922 -2976 6956
rect -3134 6916 -2976 6922
rect -2798 6956 -2640 6972
rect -2798 6922 -2783 6956
rect -2749 6922 -2689 6956
rect -2655 6922 -2640 6956
rect -2798 6916 -2640 6922
rect -5242 6326 -5226 6616
rect -5002 6326 -4984 6616
rect -5242 5762 -4984 6326
rect -4622 6872 -4470 6884
rect -4622 5896 -4584 6872
rect -4550 5896 -4510 6872
rect -4476 5896 -4470 6872
rect -4622 5884 -4470 5896
rect -4428 6874 -4370 6886
rect -4428 5896 -4416 5898
rect -4382 5896 -4370 5898
rect -4428 5884 -4370 5896
rect -4328 6872 -4134 6884
rect -4328 5896 -4322 6872
rect -4288 5896 -4248 6872
rect -4214 5896 -4174 6872
rect -4140 5896 -4134 6872
rect -4328 5884 -4134 5896
rect -4092 6874 -4034 6886
rect -4092 5896 -4080 5898
rect -4046 5896 -4034 5898
rect -4092 5884 -4034 5896
rect -3992 6872 -3798 6884
rect -3992 5896 -3986 6872
rect -3952 5896 -3912 6872
rect -3878 5896 -3838 6872
rect -3804 5896 -3798 6872
rect -3992 5884 -3798 5896
rect -3756 6874 -3698 6886
rect -3756 5896 -3744 5898
rect -3710 5896 -3698 5898
rect -3756 5884 -3698 5896
rect -3656 6872 -3462 6884
rect -3656 5896 -3650 6872
rect -3616 5896 -3576 6872
rect -3542 5896 -3502 6872
rect -3468 5896 -3462 6872
rect -3656 5884 -3462 5896
rect -3420 6874 -3362 6886
rect -3420 5896 -3408 5898
rect -3374 5896 -3362 5898
rect -3420 5884 -3362 5896
rect -3320 6872 -3126 6884
rect -3320 5896 -3314 6872
rect -3280 5896 -3240 6872
rect -3206 5896 -3166 6872
rect -3132 5896 -3126 6872
rect -3320 5884 -3126 5896
rect -3084 6874 -3026 6886
rect -3084 5896 -3072 5898
rect -3038 5896 -3026 5898
rect -3084 5884 -3026 5896
rect -2984 6872 -2790 6884
rect -2984 5896 -2978 6872
rect -2944 5896 -2904 6872
rect -2870 5896 -2830 6872
rect -2796 5896 -2790 6872
rect -2984 5884 -2790 5896
rect -2748 6874 -2690 6886
rect -2610 6884 -2498 6886
rect -2748 5896 -2736 5898
rect -2702 5896 -2690 5898
rect -2748 5884 -2690 5896
rect -2648 6872 -2498 6884
rect -2648 5896 -2642 6872
rect -2608 5896 -2568 6872
rect -2534 5896 -2498 6872
rect -2648 5884 -2498 5896
rect -4622 5762 -4510 5884
rect -4478 5846 -4320 5852
rect -4478 5812 -4463 5846
rect -4429 5812 -4369 5846
rect -4335 5812 -4320 5846
rect -4478 5806 -4320 5812
rect -4288 5762 -4176 5884
rect -4142 5846 -3984 5852
rect -4142 5812 -4127 5846
rect -4093 5812 -4033 5846
rect -3999 5812 -3984 5846
rect -4142 5806 -3984 5812
rect -3952 5762 -3840 5884
rect -3806 5846 -3648 5852
rect -3806 5812 -3791 5846
rect -3757 5812 -3697 5846
rect -3663 5812 -3648 5846
rect -3806 5806 -3648 5812
rect -3616 5762 -3504 5884
rect -3470 5846 -3312 5852
rect -3470 5812 -3455 5846
rect -3421 5812 -3361 5846
rect -3327 5812 -3312 5846
rect -3470 5806 -3312 5812
rect -3280 5762 -3168 5884
rect -3134 5846 -2976 5852
rect -3134 5812 -3119 5846
rect -3085 5812 -3025 5846
rect -2991 5812 -2976 5846
rect -3134 5806 -2976 5812
rect -2944 5762 -2832 5884
rect -2798 5846 -2640 5852
rect -2798 5812 -2783 5846
rect -2749 5812 -2689 5846
rect -2655 5812 -2640 5846
rect -2798 5806 -2640 5812
rect -2610 5762 -2498 5884
rect -5242 5756 -2498 5762
rect -5242 5704 -5200 5756
rect -2518 5704 -2498 5756
rect -5242 5698 -2498 5704
rect -5242 5674 -4984 5698
rect -2418 5612 -2306 7160
rect 450 7122 562 8704
rect 6820 8872 6932 8882
rect 6820 8704 6850 8872
rect 6906 8704 6932 8872
rect 590 8602 3086 8608
rect 590 8550 610 8602
rect 3066 8550 3086 8602
rect 590 8544 3086 8550
rect 590 8410 702 8544
rect 974 8410 1086 8544
rect 1378 8410 1490 8544
rect 1782 8410 1894 8544
rect 2186 8410 2298 8544
rect 2590 8410 2702 8544
rect 2974 8410 3086 8544
rect 590 8398 724 8410
rect 806 8408 852 8410
rect 590 7422 610 8398
rect 644 7422 684 8398
rect 718 7422 724 8398
rect 590 7410 724 7422
rect 800 8398 858 8408
rect 800 7416 858 7422
rect 934 8398 1128 8410
rect 1210 8408 1256 8410
rect 934 7422 940 8398
rect 974 7422 1014 8398
rect 1048 7422 1088 8398
rect 1122 7422 1128 8398
rect 806 7410 852 7416
rect 934 7410 1128 7422
rect 1204 8398 1262 8408
rect 1204 7416 1262 7422
rect 1338 8398 1532 8410
rect 1614 8408 1660 8410
rect 1338 7422 1344 8398
rect 1378 7422 1418 8398
rect 1452 7422 1492 8398
rect 1526 7422 1532 8398
rect 1210 7410 1256 7416
rect 1338 7410 1532 7422
rect 1608 8398 1666 8408
rect 1608 7416 1666 7422
rect 1742 8398 1936 8410
rect 2018 8408 2064 8410
rect 1742 7422 1748 8398
rect 1782 7422 1822 8398
rect 1856 7422 1896 8398
rect 1930 7422 1936 8398
rect 1614 7410 1660 7416
rect 1742 7410 1936 7422
rect 2012 8398 2070 8408
rect 2012 7416 2070 7422
rect 2146 8398 2340 8410
rect 2422 8408 2468 8410
rect 2146 7422 2152 8398
rect 2186 7422 2226 8398
rect 2260 7422 2300 8398
rect 2334 7422 2340 8398
rect 2018 7410 2064 7416
rect 2146 7410 2340 7422
rect 2416 8398 2474 8408
rect 2416 7416 2474 7422
rect 2550 8398 2744 8410
rect 2826 8408 2872 8410
rect 2550 7422 2556 8398
rect 2590 7422 2630 8398
rect 2664 7422 2704 8398
rect 2738 7422 2744 8398
rect 2422 7410 2468 7416
rect 2550 7410 2744 7422
rect 2820 8398 2878 8408
rect 2820 7416 2878 7422
rect 2954 8398 3086 8410
rect 2954 7422 2960 8398
rect 2994 7422 3034 8398
rect 3068 7422 3086 8398
rect 2826 7410 2872 7416
rect 2954 7410 3086 7422
rect 732 7363 926 7370
rect 732 7329 746 7363
rect 784 7329 874 7363
rect 912 7329 926 7363
rect 732 7310 926 7329
rect 1136 7363 1330 7370
rect 1136 7329 1150 7363
rect 1188 7329 1278 7363
rect 1316 7329 1330 7363
rect 1136 7310 1330 7329
rect 1540 7363 1734 7370
rect 1540 7329 1554 7363
rect 1592 7329 1682 7363
rect 1720 7329 1734 7363
rect 804 7268 926 7310
rect 804 7262 1054 7268
rect 1028 7210 1054 7262
rect 804 7204 1054 7210
rect 450 7064 562 7070
rect 920 7022 1054 7204
rect 1166 7128 1300 7310
rect 1540 7268 1734 7329
rect 1944 7363 2138 7370
rect 1944 7329 1958 7363
rect 1996 7329 2086 7363
rect 2124 7329 2138 7363
rect 1540 7262 1764 7268
rect 1540 7204 1764 7210
rect 1166 7122 1414 7128
rect 1390 7070 1414 7122
rect 1166 7064 1414 7070
rect 920 7006 1078 7022
rect 920 6972 935 7006
rect 969 6972 1029 7006
rect 1063 6972 1078 7006
rect 920 6966 1078 6972
rect 1256 7006 1414 7064
rect 1256 6972 1271 7006
rect 1305 6972 1365 7006
rect 1399 6972 1414 7006
rect 1256 6966 1414 6972
rect 1592 7006 1750 7204
rect 1944 7128 2138 7329
rect 2348 7363 2542 7370
rect 2348 7329 2362 7363
rect 2400 7329 2490 7363
rect 2528 7329 2542 7363
rect 2348 7268 2542 7329
rect 2294 7262 2542 7268
rect 2518 7210 2542 7262
rect 2294 7204 2542 7210
rect 2752 7363 2946 7370
rect 2752 7329 2766 7363
rect 2804 7329 2894 7363
rect 2932 7329 2946 7363
rect 2752 7292 2946 7329
rect 1920 7122 2144 7128
rect 1920 7064 2144 7070
rect 1592 6972 1607 7006
rect 1641 6972 1701 7006
rect 1735 6972 1750 7006
rect 1592 6966 1750 6972
rect 1928 7006 2086 7064
rect 2294 7022 2406 7204
rect 2752 7128 2872 7292
rect 2640 7122 2872 7128
rect 2864 7070 2872 7122
rect 2640 7064 2872 7070
rect 2980 7262 3092 7268
rect 2640 7022 2758 7064
rect 1928 6972 1943 7006
rect 1977 6972 2037 7006
rect 2071 6972 2086 7006
rect 1928 6966 2086 6972
rect 2264 7006 2422 7022
rect 2264 6972 2279 7006
rect 2313 6972 2373 7006
rect 2407 6972 2422 7006
rect 2264 6966 2422 6972
rect 2600 7006 2758 7022
rect 2600 6972 2615 7006
rect 2649 6972 2709 7006
rect 2743 6972 2758 7006
rect 2600 6966 2758 6972
rect -1684 6614 -1180 6664
rect -1684 6324 -1422 6614
rect -1198 6324 -1180 6614
rect -1684 5806 -1180 6324
rect 792 6642 848 6934
rect 876 6928 934 6934
rect 876 6664 888 6670
rect 792 6634 854 6642
rect 792 5946 814 6634
rect 848 5946 854 6634
rect 792 5812 854 5946
rect 882 5946 888 6664
rect 922 6664 934 6670
rect 976 6922 1022 6934
rect 922 5946 928 6664
rect 976 6330 982 6922
rect 882 5934 928 5946
rect 970 6320 982 6330
rect 1016 6330 1022 6922
rect 1064 6928 1122 6934
rect 1064 6664 1076 6670
rect 1016 6320 1028 6330
rect 970 5946 982 5948
rect 1016 5946 1028 5948
rect 970 5934 1028 5946
rect 1070 5946 1076 6664
rect 1110 6664 1122 6670
rect 1110 5946 1116 6664
rect 1150 6640 1184 6934
rect 1212 6928 1270 6934
rect 1212 6664 1224 6670
rect 1070 5934 1116 5946
rect 1144 6634 1190 6640
rect 1144 5946 1150 6634
rect 1184 5946 1190 6634
rect 1144 5812 1190 5946
rect 1218 5946 1224 6664
rect 1258 6664 1270 6670
rect 1312 6922 1358 6934
rect 1258 5946 1264 6664
rect 1312 6330 1318 6922
rect 1218 5934 1264 5946
rect 1306 6320 1318 6330
rect 1352 6330 1358 6922
rect 1400 6928 1458 6934
rect 1400 6664 1412 6670
rect 1352 6320 1364 6330
rect 1306 5946 1318 5948
rect 1352 5946 1364 5948
rect 1306 5934 1364 5946
rect 1406 5946 1412 6664
rect 1446 6664 1458 6670
rect 1446 5946 1452 6664
rect 1486 6640 1520 6934
rect 1548 6928 1606 6934
rect 1548 6664 1560 6670
rect 1406 5934 1452 5946
rect 1480 6634 1526 6640
rect 1480 5946 1486 6634
rect 1520 5946 1526 6634
rect 1480 5812 1526 5946
rect 1554 5946 1560 6664
rect 1594 6664 1606 6670
rect 1648 6922 1694 6934
rect 1594 5946 1600 6664
rect 1648 6330 1654 6922
rect 1554 5934 1600 5946
rect 1642 6320 1654 6330
rect 1688 6330 1694 6922
rect 1736 6928 1794 6934
rect 1736 6664 1748 6670
rect 1688 6320 1700 6330
rect 1642 5946 1654 5948
rect 1688 5946 1700 5948
rect 1642 5934 1700 5946
rect 1742 5946 1748 6664
rect 1782 6664 1794 6670
rect 1782 5946 1788 6664
rect 1822 6640 1856 6934
rect 1884 6928 1942 6934
rect 1884 6664 1896 6670
rect 1742 5934 1788 5946
rect 1816 6634 1862 6640
rect 1816 5946 1822 6634
rect 1856 5946 1862 6634
rect 1816 5812 1862 5946
rect 1890 5946 1896 6664
rect 1930 6664 1942 6670
rect 1984 6922 2030 6934
rect 1930 5946 1936 6664
rect 1984 6330 1990 6922
rect 1890 5934 1936 5946
rect 1978 6320 1990 6330
rect 2024 6330 2030 6922
rect 2072 6928 2130 6934
rect 2072 6664 2084 6670
rect 2024 6320 2036 6330
rect 1978 5946 1990 5948
rect 2024 5946 2036 5948
rect 1978 5934 2036 5946
rect 2078 5946 2084 6664
rect 2118 6664 2130 6670
rect 2118 5946 2124 6664
rect 2158 6640 2192 6934
rect 2220 6928 2278 6934
rect 2220 6664 2232 6670
rect 2078 5934 2124 5946
rect 2152 6634 2198 6640
rect 2152 5946 2158 6634
rect 2192 5946 2198 6634
rect 2152 5812 2198 5946
rect 2226 5946 2232 6664
rect 2266 6664 2278 6670
rect 2320 6922 2366 6934
rect 2266 5946 2272 6664
rect 2320 6330 2326 6922
rect 2226 5934 2272 5946
rect 2314 6320 2326 6330
rect 2360 6330 2366 6922
rect 2408 6928 2466 6934
rect 2408 6664 2420 6670
rect 2360 6320 2372 6330
rect 2314 5946 2326 5948
rect 2360 5946 2372 5948
rect 2314 5934 2372 5946
rect 2414 5946 2420 6664
rect 2454 6664 2466 6670
rect 2454 5946 2460 6664
rect 2494 6640 2528 6934
rect 2556 6928 2614 6934
rect 2556 6664 2568 6670
rect 2414 5934 2460 5946
rect 2488 6634 2534 6640
rect 2488 5946 2494 6634
rect 2528 5946 2534 6634
rect 2488 5812 2534 5946
rect 2562 5946 2568 6664
rect 2602 6664 2614 6670
rect 2656 6922 2702 6934
rect 2602 5946 2608 6664
rect 2656 6330 2662 6922
rect 2562 5934 2608 5946
rect 2650 6320 2662 6330
rect 2696 6330 2702 6922
rect 2744 6928 2802 6934
rect 2744 6664 2756 6670
rect 2696 6320 2708 6330
rect 2650 5946 2662 5948
rect 2696 5946 2708 5948
rect 2650 5934 2708 5946
rect 2750 5946 2756 6664
rect 2790 6664 2802 6670
rect 2790 5946 2796 6664
rect 2830 6640 2886 6934
rect 2750 5934 2796 5946
rect 2824 6634 2886 6640
rect 2824 5946 2830 6634
rect 2864 5946 2886 6634
rect 2824 5812 2886 5946
rect -1684 5754 -1656 5806
rect -1208 5754 -1180 5806
rect -1684 5724 -1180 5754
rect 776 5806 2900 5812
rect 776 5754 796 5806
rect 2880 5754 2900 5806
rect 776 5748 2900 5754
rect -2418 5444 -2390 5612
rect -2334 5444 -2306 5612
rect 2980 5662 3092 7210
rect 6820 7122 6932 8704
rect 13190 8872 13302 8882
rect 13190 8704 13220 8872
rect 13276 8704 13302 8872
rect 6960 8602 9456 8608
rect 6960 8550 6980 8602
rect 9436 8550 9456 8602
rect 6960 8544 9456 8550
rect 6960 8410 7072 8544
rect 7344 8410 7456 8544
rect 7748 8410 7860 8544
rect 8152 8410 8264 8544
rect 8556 8410 8668 8544
rect 8960 8410 9072 8544
rect 9344 8410 9456 8544
rect 6960 8398 7094 8410
rect 7176 8408 7222 8410
rect 6960 7422 6980 8398
rect 7014 7422 7054 8398
rect 7088 7422 7094 8398
rect 6960 7410 7094 7422
rect 7170 8398 7228 8408
rect 7170 7416 7228 7422
rect 7304 8398 7498 8410
rect 7580 8408 7626 8410
rect 7304 7422 7310 8398
rect 7344 7422 7384 8398
rect 7418 7422 7458 8398
rect 7492 7422 7498 8398
rect 7176 7410 7222 7416
rect 7304 7410 7498 7422
rect 7574 8398 7632 8408
rect 7574 7416 7632 7422
rect 7708 8398 7902 8410
rect 7984 8408 8030 8410
rect 7708 7422 7714 8398
rect 7748 7422 7788 8398
rect 7822 7422 7862 8398
rect 7896 7422 7902 8398
rect 7580 7410 7626 7416
rect 7708 7410 7902 7422
rect 7978 8398 8036 8408
rect 7978 7416 8036 7422
rect 8112 8398 8306 8410
rect 8388 8408 8434 8410
rect 8112 7422 8118 8398
rect 8152 7422 8192 8398
rect 8226 7422 8266 8398
rect 8300 7422 8306 8398
rect 7984 7410 8030 7416
rect 8112 7410 8306 7422
rect 8382 8398 8440 8408
rect 8382 7416 8440 7422
rect 8516 8398 8710 8410
rect 8792 8408 8838 8410
rect 8516 7422 8522 8398
rect 8556 7422 8596 8398
rect 8630 7422 8670 8398
rect 8704 7422 8710 8398
rect 8388 7410 8434 7416
rect 8516 7410 8710 7422
rect 8786 8398 8844 8408
rect 8786 7416 8844 7422
rect 8920 8398 9114 8410
rect 9196 8408 9242 8410
rect 8920 7422 8926 8398
rect 8960 7422 9000 8398
rect 9034 7422 9074 8398
rect 9108 7422 9114 8398
rect 8792 7410 8838 7416
rect 8920 7410 9114 7422
rect 9190 8398 9248 8408
rect 9190 7416 9248 7422
rect 9324 8398 9456 8410
rect 9324 7422 9330 8398
rect 9364 7422 9404 8398
rect 9438 7422 9456 8398
rect 9196 7410 9242 7416
rect 9324 7410 9456 7422
rect 7102 7363 7296 7370
rect 7102 7329 7116 7363
rect 7154 7329 7244 7363
rect 7282 7329 7296 7363
rect 7102 7310 7296 7329
rect 7506 7363 7700 7370
rect 7506 7329 7520 7363
rect 7558 7329 7648 7363
rect 7686 7329 7700 7363
rect 7506 7310 7700 7329
rect 7910 7363 8104 7370
rect 7910 7329 7924 7363
rect 7962 7329 8052 7363
rect 8090 7329 8104 7363
rect 7174 7268 7296 7310
rect 7174 7262 7424 7268
rect 7398 7210 7424 7262
rect 7174 7204 7424 7210
rect 6820 7064 6932 7070
rect 7290 7022 7424 7204
rect 7536 7128 7670 7310
rect 7910 7268 8104 7329
rect 8314 7363 8508 7370
rect 8314 7329 8328 7363
rect 8366 7329 8456 7363
rect 8494 7329 8508 7363
rect 7910 7262 8134 7268
rect 7910 7204 8134 7210
rect 7536 7122 7784 7128
rect 7760 7070 7784 7122
rect 7536 7064 7784 7070
rect 7290 7006 7448 7022
rect 7290 6972 7305 7006
rect 7339 6972 7399 7006
rect 7433 6972 7448 7006
rect 7290 6966 7448 6972
rect 7626 7006 7784 7064
rect 7626 6972 7641 7006
rect 7675 6972 7735 7006
rect 7769 6972 7784 7006
rect 7626 6966 7784 6972
rect 7962 7006 8120 7204
rect 8314 7128 8508 7329
rect 8718 7363 8912 7370
rect 8718 7329 8732 7363
rect 8770 7329 8860 7363
rect 8898 7329 8912 7363
rect 8718 7268 8912 7329
rect 8664 7262 8912 7268
rect 8888 7210 8912 7262
rect 8664 7204 8912 7210
rect 9122 7363 9316 7370
rect 9122 7329 9136 7363
rect 9174 7329 9264 7363
rect 9302 7329 9316 7363
rect 9122 7292 9316 7329
rect 8290 7122 8514 7128
rect 8290 7064 8514 7070
rect 7962 6972 7977 7006
rect 8011 6972 8071 7006
rect 8105 6972 8120 7006
rect 7962 6966 8120 6972
rect 8298 7006 8456 7064
rect 8664 7022 8776 7204
rect 9122 7128 9242 7292
rect 9010 7122 9242 7128
rect 9234 7070 9242 7122
rect 9010 7064 9242 7070
rect 9350 7262 9462 7268
rect 9010 7022 9128 7064
rect 8298 6972 8313 7006
rect 8347 6972 8407 7006
rect 8441 6972 8456 7006
rect 8298 6966 8456 6972
rect 8634 7006 8792 7022
rect 8634 6972 8649 7006
rect 8683 6972 8743 7006
rect 8777 6972 8792 7006
rect 8634 6966 8792 6972
rect 8970 7006 9128 7022
rect 8970 6972 8985 7006
rect 9019 6972 9079 7006
rect 9113 6972 9128 7006
rect 8970 6966 9128 6972
rect 4686 6614 5190 6664
rect 4686 6324 4948 6614
rect 5172 6324 5190 6614
rect 4686 5806 5190 6324
rect 7162 6642 7218 6934
rect 7246 6928 7304 6934
rect 7246 6664 7258 6670
rect 7162 6634 7224 6642
rect 7162 5946 7184 6634
rect 7218 5946 7224 6634
rect 7162 5812 7224 5946
rect 7252 5946 7258 6664
rect 7292 6664 7304 6670
rect 7346 6922 7392 6934
rect 7292 5946 7298 6664
rect 7346 6330 7352 6922
rect 7252 5934 7298 5946
rect 7340 6320 7352 6330
rect 7386 6330 7392 6922
rect 7434 6928 7492 6934
rect 7434 6664 7446 6670
rect 7386 6320 7398 6330
rect 7340 5946 7352 5948
rect 7386 5946 7398 5948
rect 7340 5934 7398 5946
rect 7440 5946 7446 6664
rect 7480 6664 7492 6670
rect 7480 5946 7486 6664
rect 7520 6640 7554 6934
rect 7582 6928 7640 6934
rect 7582 6664 7594 6670
rect 7440 5934 7486 5946
rect 7514 6634 7560 6640
rect 7514 5946 7520 6634
rect 7554 5946 7560 6634
rect 7514 5812 7560 5946
rect 7588 5946 7594 6664
rect 7628 6664 7640 6670
rect 7682 6922 7728 6934
rect 7628 5946 7634 6664
rect 7682 6330 7688 6922
rect 7588 5934 7634 5946
rect 7676 6320 7688 6330
rect 7722 6330 7728 6922
rect 7770 6928 7828 6934
rect 7770 6664 7782 6670
rect 7722 6320 7734 6330
rect 7676 5946 7688 5948
rect 7722 5946 7734 5948
rect 7676 5934 7734 5946
rect 7776 5946 7782 6664
rect 7816 6664 7828 6670
rect 7816 5946 7822 6664
rect 7856 6640 7890 6934
rect 7918 6928 7976 6934
rect 7918 6664 7930 6670
rect 7776 5934 7822 5946
rect 7850 6634 7896 6640
rect 7850 5946 7856 6634
rect 7890 5946 7896 6634
rect 7850 5812 7896 5946
rect 7924 5946 7930 6664
rect 7964 6664 7976 6670
rect 8018 6922 8064 6934
rect 7964 5946 7970 6664
rect 8018 6330 8024 6922
rect 7924 5934 7970 5946
rect 8012 6320 8024 6330
rect 8058 6330 8064 6922
rect 8106 6928 8164 6934
rect 8106 6664 8118 6670
rect 8058 6320 8070 6330
rect 8012 5946 8024 5948
rect 8058 5946 8070 5948
rect 8012 5934 8070 5946
rect 8112 5946 8118 6664
rect 8152 6664 8164 6670
rect 8152 5946 8158 6664
rect 8192 6640 8226 6934
rect 8254 6928 8312 6934
rect 8254 6664 8266 6670
rect 8112 5934 8158 5946
rect 8186 6634 8232 6640
rect 8186 5946 8192 6634
rect 8226 5946 8232 6634
rect 8186 5812 8232 5946
rect 8260 5946 8266 6664
rect 8300 6664 8312 6670
rect 8354 6922 8400 6934
rect 8300 5946 8306 6664
rect 8354 6330 8360 6922
rect 8260 5934 8306 5946
rect 8348 6320 8360 6330
rect 8394 6330 8400 6922
rect 8442 6928 8500 6934
rect 8442 6664 8454 6670
rect 8394 6320 8406 6330
rect 8348 5946 8360 5948
rect 8394 5946 8406 5948
rect 8348 5934 8406 5946
rect 8448 5946 8454 6664
rect 8488 6664 8500 6670
rect 8488 5946 8494 6664
rect 8528 6640 8562 6934
rect 8590 6928 8648 6934
rect 8590 6664 8602 6670
rect 8448 5934 8494 5946
rect 8522 6634 8568 6640
rect 8522 5946 8528 6634
rect 8562 5946 8568 6634
rect 8522 5812 8568 5946
rect 8596 5946 8602 6664
rect 8636 6664 8648 6670
rect 8690 6922 8736 6934
rect 8636 5946 8642 6664
rect 8690 6330 8696 6922
rect 8596 5934 8642 5946
rect 8684 6320 8696 6330
rect 8730 6330 8736 6922
rect 8778 6928 8836 6934
rect 8778 6664 8790 6670
rect 8730 6320 8742 6330
rect 8684 5946 8696 5948
rect 8730 5946 8742 5948
rect 8684 5934 8742 5946
rect 8784 5946 8790 6664
rect 8824 6664 8836 6670
rect 8824 5946 8830 6664
rect 8864 6640 8898 6934
rect 8926 6928 8984 6934
rect 8926 6664 8938 6670
rect 8784 5934 8830 5946
rect 8858 6634 8904 6640
rect 8858 5946 8864 6634
rect 8898 5946 8904 6634
rect 8858 5812 8904 5946
rect 8932 5946 8938 6664
rect 8972 6664 8984 6670
rect 9026 6922 9072 6934
rect 8972 5946 8978 6664
rect 9026 6330 9032 6922
rect 8932 5934 8978 5946
rect 9020 6320 9032 6330
rect 9066 6330 9072 6922
rect 9114 6928 9172 6934
rect 9114 6664 9126 6670
rect 9066 6320 9078 6330
rect 9020 5946 9032 5948
rect 9066 5946 9078 5948
rect 9020 5934 9078 5946
rect 9120 5946 9126 6664
rect 9160 6664 9172 6670
rect 9160 5946 9166 6664
rect 9200 6640 9256 6934
rect 9120 5934 9166 5946
rect 9194 6634 9256 6640
rect 9194 5946 9200 6634
rect 9234 5946 9256 6634
rect 9194 5812 9256 5946
rect 4686 5754 4714 5806
rect 5162 5754 5190 5806
rect 4686 5724 5190 5754
rect 7146 5806 9270 5812
rect 7146 5754 7166 5806
rect 9250 5754 9270 5806
rect 7146 5748 9270 5754
rect 2980 5494 3008 5662
rect 3064 5494 3092 5662
rect 2980 5484 3092 5494
rect 9350 5662 9462 7210
rect 13190 7122 13302 8704
rect 19560 8872 19672 8882
rect 19560 8704 19590 8872
rect 19646 8704 19672 8872
rect 13330 8602 15826 8608
rect 13330 8550 13350 8602
rect 15806 8550 15826 8602
rect 13330 8544 15826 8550
rect 13330 8410 13442 8544
rect 13714 8410 13826 8544
rect 14118 8410 14230 8544
rect 14522 8410 14634 8544
rect 14926 8410 15038 8544
rect 15330 8410 15442 8544
rect 15714 8410 15826 8544
rect 13330 8398 13464 8410
rect 13546 8408 13592 8410
rect 13330 7422 13350 8398
rect 13384 7422 13424 8398
rect 13458 7422 13464 8398
rect 13330 7410 13464 7422
rect 13540 8398 13598 8408
rect 13540 7416 13598 7422
rect 13674 8398 13868 8410
rect 13950 8408 13996 8410
rect 13674 7422 13680 8398
rect 13714 7422 13754 8398
rect 13788 7422 13828 8398
rect 13862 7422 13868 8398
rect 13546 7410 13592 7416
rect 13674 7410 13868 7422
rect 13944 8398 14002 8408
rect 13944 7416 14002 7422
rect 14078 8398 14272 8410
rect 14354 8408 14400 8410
rect 14078 7422 14084 8398
rect 14118 7422 14158 8398
rect 14192 7422 14232 8398
rect 14266 7422 14272 8398
rect 13950 7410 13996 7416
rect 14078 7410 14272 7422
rect 14348 8398 14406 8408
rect 14348 7416 14406 7422
rect 14482 8398 14676 8410
rect 14758 8408 14804 8410
rect 14482 7422 14488 8398
rect 14522 7422 14562 8398
rect 14596 7422 14636 8398
rect 14670 7422 14676 8398
rect 14354 7410 14400 7416
rect 14482 7410 14676 7422
rect 14752 8398 14810 8408
rect 14752 7416 14810 7422
rect 14886 8398 15080 8410
rect 15162 8408 15208 8410
rect 14886 7422 14892 8398
rect 14926 7422 14966 8398
rect 15000 7422 15040 8398
rect 15074 7422 15080 8398
rect 14758 7410 14804 7416
rect 14886 7410 15080 7422
rect 15156 8398 15214 8408
rect 15156 7416 15214 7422
rect 15290 8398 15484 8410
rect 15566 8408 15612 8410
rect 15290 7422 15296 8398
rect 15330 7422 15370 8398
rect 15404 7422 15444 8398
rect 15478 7422 15484 8398
rect 15162 7410 15208 7416
rect 15290 7410 15484 7422
rect 15560 8398 15618 8408
rect 15560 7416 15618 7422
rect 15694 8398 15826 8410
rect 15694 7422 15700 8398
rect 15734 7422 15774 8398
rect 15808 7422 15826 8398
rect 15566 7410 15612 7416
rect 15694 7410 15826 7422
rect 13472 7363 13666 7370
rect 13472 7329 13486 7363
rect 13524 7329 13614 7363
rect 13652 7329 13666 7363
rect 13472 7310 13666 7329
rect 13876 7363 14070 7370
rect 13876 7329 13890 7363
rect 13928 7329 14018 7363
rect 14056 7329 14070 7363
rect 13876 7310 14070 7329
rect 14280 7363 14474 7370
rect 14280 7329 14294 7363
rect 14332 7329 14422 7363
rect 14460 7329 14474 7363
rect 13544 7268 13666 7310
rect 13544 7262 13794 7268
rect 13768 7210 13794 7262
rect 13544 7204 13794 7210
rect 13190 7064 13302 7070
rect 13660 7022 13794 7204
rect 13906 7128 14040 7310
rect 14280 7268 14474 7329
rect 14684 7363 14878 7370
rect 14684 7329 14698 7363
rect 14736 7329 14826 7363
rect 14864 7329 14878 7363
rect 14280 7262 14504 7268
rect 14280 7204 14504 7210
rect 13906 7122 14154 7128
rect 14130 7070 14154 7122
rect 13906 7064 14154 7070
rect 13660 7006 13818 7022
rect 13660 6972 13675 7006
rect 13709 6972 13769 7006
rect 13803 6972 13818 7006
rect 13660 6966 13818 6972
rect 13996 7006 14154 7064
rect 13996 6972 14011 7006
rect 14045 6972 14105 7006
rect 14139 6972 14154 7006
rect 13996 6966 14154 6972
rect 14332 7006 14490 7204
rect 14684 7128 14878 7329
rect 15088 7363 15282 7370
rect 15088 7329 15102 7363
rect 15140 7329 15230 7363
rect 15268 7329 15282 7363
rect 15088 7268 15282 7329
rect 15034 7262 15282 7268
rect 15258 7210 15282 7262
rect 15034 7204 15282 7210
rect 15492 7363 15686 7370
rect 15492 7329 15506 7363
rect 15544 7329 15634 7363
rect 15672 7329 15686 7363
rect 15492 7292 15686 7329
rect 14660 7122 14884 7128
rect 14660 7064 14884 7070
rect 14332 6972 14347 7006
rect 14381 6972 14441 7006
rect 14475 6972 14490 7006
rect 14332 6966 14490 6972
rect 14668 7006 14826 7064
rect 15034 7022 15146 7204
rect 15492 7128 15612 7292
rect 15380 7122 15612 7128
rect 15604 7070 15612 7122
rect 15380 7064 15612 7070
rect 15720 7262 15832 7268
rect 15380 7022 15498 7064
rect 14668 6972 14683 7006
rect 14717 6972 14777 7006
rect 14811 6972 14826 7006
rect 14668 6966 14826 6972
rect 15004 7006 15162 7022
rect 15004 6972 15019 7006
rect 15053 6972 15113 7006
rect 15147 6972 15162 7006
rect 15004 6966 15162 6972
rect 15340 7006 15498 7022
rect 15340 6972 15355 7006
rect 15389 6972 15449 7006
rect 15483 6972 15498 7006
rect 15340 6966 15498 6972
rect 11056 6614 11560 6664
rect 11056 6324 11318 6614
rect 11542 6324 11560 6614
rect 11056 5806 11560 6324
rect 13532 6642 13588 6934
rect 13616 6928 13674 6934
rect 13616 6664 13628 6670
rect 13532 6634 13594 6642
rect 13532 5946 13554 6634
rect 13588 5946 13594 6634
rect 13532 5812 13594 5946
rect 13622 5946 13628 6664
rect 13662 6664 13674 6670
rect 13716 6922 13762 6934
rect 13662 5946 13668 6664
rect 13716 6330 13722 6922
rect 13622 5934 13668 5946
rect 13710 6320 13722 6330
rect 13756 6330 13762 6922
rect 13804 6928 13862 6934
rect 13804 6664 13816 6670
rect 13756 6320 13768 6330
rect 13710 5946 13722 5948
rect 13756 5946 13768 5948
rect 13710 5934 13768 5946
rect 13810 5946 13816 6664
rect 13850 6664 13862 6670
rect 13850 5946 13856 6664
rect 13890 6640 13924 6934
rect 13952 6928 14010 6934
rect 13952 6664 13964 6670
rect 13810 5934 13856 5946
rect 13884 6634 13930 6640
rect 13884 5946 13890 6634
rect 13924 5946 13930 6634
rect 13884 5812 13930 5946
rect 13958 5946 13964 6664
rect 13998 6664 14010 6670
rect 14052 6922 14098 6934
rect 13998 5946 14004 6664
rect 14052 6330 14058 6922
rect 13958 5934 14004 5946
rect 14046 6320 14058 6330
rect 14092 6330 14098 6922
rect 14140 6928 14198 6934
rect 14140 6664 14152 6670
rect 14092 6320 14104 6330
rect 14046 5946 14058 5948
rect 14092 5946 14104 5948
rect 14046 5934 14104 5946
rect 14146 5946 14152 6664
rect 14186 6664 14198 6670
rect 14186 5946 14192 6664
rect 14226 6640 14260 6934
rect 14288 6928 14346 6934
rect 14288 6664 14300 6670
rect 14146 5934 14192 5946
rect 14220 6634 14266 6640
rect 14220 5946 14226 6634
rect 14260 5946 14266 6634
rect 14220 5812 14266 5946
rect 14294 5946 14300 6664
rect 14334 6664 14346 6670
rect 14388 6922 14434 6934
rect 14334 5946 14340 6664
rect 14388 6330 14394 6922
rect 14294 5934 14340 5946
rect 14382 6320 14394 6330
rect 14428 6330 14434 6922
rect 14476 6928 14534 6934
rect 14476 6664 14488 6670
rect 14428 6320 14440 6330
rect 14382 5946 14394 5948
rect 14428 5946 14440 5948
rect 14382 5934 14440 5946
rect 14482 5946 14488 6664
rect 14522 6664 14534 6670
rect 14522 5946 14528 6664
rect 14562 6640 14596 6934
rect 14624 6928 14682 6934
rect 14624 6664 14636 6670
rect 14482 5934 14528 5946
rect 14556 6634 14602 6640
rect 14556 5946 14562 6634
rect 14596 5946 14602 6634
rect 14556 5812 14602 5946
rect 14630 5946 14636 6664
rect 14670 6664 14682 6670
rect 14724 6922 14770 6934
rect 14670 5946 14676 6664
rect 14724 6330 14730 6922
rect 14630 5934 14676 5946
rect 14718 6320 14730 6330
rect 14764 6330 14770 6922
rect 14812 6928 14870 6934
rect 14812 6664 14824 6670
rect 14764 6320 14776 6330
rect 14718 5946 14730 5948
rect 14764 5946 14776 5948
rect 14718 5934 14776 5946
rect 14818 5946 14824 6664
rect 14858 6664 14870 6670
rect 14858 5946 14864 6664
rect 14898 6640 14932 6934
rect 14960 6928 15018 6934
rect 14960 6664 14972 6670
rect 14818 5934 14864 5946
rect 14892 6634 14938 6640
rect 14892 5946 14898 6634
rect 14932 5946 14938 6634
rect 14892 5812 14938 5946
rect 14966 5946 14972 6664
rect 15006 6664 15018 6670
rect 15060 6922 15106 6934
rect 15006 5946 15012 6664
rect 15060 6330 15066 6922
rect 14966 5934 15012 5946
rect 15054 6320 15066 6330
rect 15100 6330 15106 6922
rect 15148 6928 15206 6934
rect 15148 6664 15160 6670
rect 15100 6320 15112 6330
rect 15054 5946 15066 5948
rect 15100 5946 15112 5948
rect 15054 5934 15112 5946
rect 15154 5946 15160 6664
rect 15194 6664 15206 6670
rect 15194 5946 15200 6664
rect 15234 6640 15268 6934
rect 15296 6928 15354 6934
rect 15296 6664 15308 6670
rect 15154 5934 15200 5946
rect 15228 6634 15274 6640
rect 15228 5946 15234 6634
rect 15268 5946 15274 6634
rect 15228 5812 15274 5946
rect 15302 5946 15308 6664
rect 15342 6664 15354 6670
rect 15396 6922 15442 6934
rect 15342 5946 15348 6664
rect 15396 6330 15402 6922
rect 15302 5934 15348 5946
rect 15390 6320 15402 6330
rect 15436 6330 15442 6922
rect 15484 6928 15542 6934
rect 15484 6664 15496 6670
rect 15436 6320 15448 6330
rect 15390 5946 15402 5948
rect 15436 5946 15448 5948
rect 15390 5934 15448 5946
rect 15490 5946 15496 6664
rect 15530 6664 15542 6670
rect 15530 5946 15536 6664
rect 15570 6640 15626 6934
rect 15490 5934 15536 5946
rect 15564 6634 15626 6640
rect 15564 5946 15570 6634
rect 15604 5946 15626 6634
rect 15564 5812 15626 5946
rect 11056 5754 11084 5806
rect 11532 5754 11560 5806
rect 11056 5724 11560 5754
rect 13516 5806 15640 5812
rect 13516 5754 13536 5806
rect 15620 5754 15640 5806
rect 13516 5748 15640 5754
rect 9350 5494 9378 5662
rect 9434 5494 9462 5662
rect 9350 5484 9462 5494
rect 15720 5662 15832 7210
rect 19560 7122 19672 8704
rect 28818 8872 28930 8882
rect 28818 8704 28848 8872
rect 28904 8704 28930 8872
rect 19700 8602 22196 8608
rect 19700 8550 19720 8602
rect 22176 8550 22196 8602
rect 19700 8544 22196 8550
rect 19700 8410 19812 8544
rect 20084 8410 20196 8544
rect 20488 8410 20600 8544
rect 20892 8410 21004 8544
rect 21296 8410 21408 8544
rect 21700 8410 21812 8544
rect 22084 8410 22196 8544
rect 19700 8398 19834 8410
rect 19916 8408 19962 8410
rect 19700 7422 19720 8398
rect 19754 7422 19794 8398
rect 19828 7422 19834 8398
rect 19700 7410 19834 7422
rect 19910 8398 19968 8408
rect 19910 7416 19968 7422
rect 20044 8398 20238 8410
rect 20320 8408 20366 8410
rect 20044 7422 20050 8398
rect 20084 7422 20124 8398
rect 20158 7422 20198 8398
rect 20232 7422 20238 8398
rect 19916 7410 19962 7416
rect 20044 7410 20238 7422
rect 20314 8398 20372 8408
rect 20314 7416 20372 7422
rect 20448 8398 20642 8410
rect 20724 8408 20770 8410
rect 20448 7422 20454 8398
rect 20488 7422 20528 8398
rect 20562 7422 20602 8398
rect 20636 7422 20642 8398
rect 20320 7410 20366 7416
rect 20448 7410 20642 7422
rect 20718 8398 20776 8408
rect 20718 7416 20776 7422
rect 20852 8398 21046 8410
rect 21128 8408 21174 8410
rect 20852 7422 20858 8398
rect 20892 7422 20932 8398
rect 20966 7422 21006 8398
rect 21040 7422 21046 8398
rect 20724 7410 20770 7416
rect 20852 7410 21046 7422
rect 21122 8398 21180 8408
rect 21122 7416 21180 7422
rect 21256 8398 21450 8410
rect 21532 8408 21578 8410
rect 21256 7422 21262 8398
rect 21296 7422 21336 8398
rect 21370 7422 21410 8398
rect 21444 7422 21450 8398
rect 21128 7410 21174 7416
rect 21256 7410 21450 7422
rect 21526 8398 21584 8408
rect 21526 7416 21584 7422
rect 21660 8398 21854 8410
rect 21936 8408 21982 8410
rect 21660 7422 21666 8398
rect 21700 7422 21740 8398
rect 21774 7422 21814 8398
rect 21848 7422 21854 8398
rect 21532 7410 21578 7416
rect 21660 7410 21854 7422
rect 21930 8398 21988 8408
rect 21930 7416 21988 7422
rect 22064 8398 22196 8410
rect 22064 7422 22070 8398
rect 22104 7422 22144 8398
rect 22178 7422 22196 8398
rect 21936 7410 21982 7416
rect 22064 7410 22196 7422
rect 19842 7363 20036 7370
rect 19842 7329 19856 7363
rect 19894 7329 19984 7363
rect 20022 7329 20036 7363
rect 19842 7310 20036 7329
rect 20246 7363 20440 7370
rect 20246 7329 20260 7363
rect 20298 7329 20388 7363
rect 20426 7329 20440 7363
rect 20246 7310 20440 7329
rect 20650 7363 20844 7370
rect 20650 7329 20664 7363
rect 20702 7329 20792 7363
rect 20830 7329 20844 7363
rect 19914 7268 20036 7310
rect 19914 7262 20164 7268
rect 20138 7210 20164 7262
rect 19914 7204 20164 7210
rect 19560 7064 19672 7070
rect 20030 7022 20164 7204
rect 20276 7128 20410 7310
rect 20650 7268 20844 7329
rect 21054 7363 21248 7370
rect 21054 7329 21068 7363
rect 21106 7329 21196 7363
rect 21234 7329 21248 7363
rect 20650 7262 20874 7268
rect 20650 7204 20874 7210
rect 20276 7122 20524 7128
rect 20500 7070 20524 7122
rect 20276 7064 20524 7070
rect 20030 7006 20188 7022
rect 20030 6972 20045 7006
rect 20079 6972 20139 7006
rect 20173 6972 20188 7006
rect 20030 6966 20188 6972
rect 20366 7006 20524 7064
rect 20366 6972 20381 7006
rect 20415 6972 20475 7006
rect 20509 6972 20524 7006
rect 20366 6966 20524 6972
rect 20702 7006 20860 7204
rect 21054 7128 21248 7329
rect 21458 7363 21652 7370
rect 21458 7329 21472 7363
rect 21510 7329 21600 7363
rect 21638 7329 21652 7363
rect 21458 7268 21652 7329
rect 21404 7262 21652 7268
rect 21628 7210 21652 7262
rect 21404 7204 21652 7210
rect 21862 7363 22056 7370
rect 21862 7329 21876 7363
rect 21914 7329 22004 7363
rect 22042 7329 22056 7363
rect 21862 7292 22056 7329
rect 21030 7122 21254 7128
rect 21030 7064 21254 7070
rect 20702 6972 20717 7006
rect 20751 6972 20811 7006
rect 20845 6972 20860 7006
rect 20702 6966 20860 6972
rect 21038 7006 21196 7064
rect 21404 7022 21516 7204
rect 21862 7128 21982 7292
rect 21750 7122 21982 7128
rect 21974 7070 21982 7122
rect 21750 7064 21982 7070
rect 22090 7262 22202 7268
rect 21750 7022 21868 7064
rect 21038 6972 21053 7006
rect 21087 6972 21147 7006
rect 21181 6972 21196 7006
rect 21038 6966 21196 6972
rect 21374 7006 21532 7022
rect 21374 6972 21389 7006
rect 21423 6972 21483 7006
rect 21517 6972 21532 7006
rect 21374 6966 21532 6972
rect 21710 7006 21868 7022
rect 21710 6972 21725 7006
rect 21759 6972 21819 7006
rect 21853 6972 21868 7006
rect 21710 6966 21868 6972
rect 17426 6614 17930 6664
rect 17426 6324 17688 6614
rect 17912 6324 17930 6614
rect 17426 5806 17930 6324
rect 19902 6642 19958 6934
rect 19986 6928 20044 6934
rect 19986 6664 19998 6670
rect 19902 6634 19964 6642
rect 19902 5946 19924 6634
rect 19958 5946 19964 6634
rect 19902 5812 19964 5946
rect 19992 5946 19998 6664
rect 20032 6664 20044 6670
rect 20086 6922 20132 6934
rect 20032 5946 20038 6664
rect 20086 6330 20092 6922
rect 19992 5934 20038 5946
rect 20080 6320 20092 6330
rect 20126 6330 20132 6922
rect 20174 6928 20232 6934
rect 20174 6664 20186 6670
rect 20126 6320 20138 6330
rect 20080 5946 20092 5948
rect 20126 5946 20138 5948
rect 20080 5934 20138 5946
rect 20180 5946 20186 6664
rect 20220 6664 20232 6670
rect 20220 5946 20226 6664
rect 20260 6640 20294 6934
rect 20322 6928 20380 6934
rect 20322 6664 20334 6670
rect 20180 5934 20226 5946
rect 20254 6634 20300 6640
rect 20254 5946 20260 6634
rect 20294 5946 20300 6634
rect 20254 5812 20300 5946
rect 20328 5946 20334 6664
rect 20368 6664 20380 6670
rect 20422 6922 20468 6934
rect 20368 5946 20374 6664
rect 20422 6330 20428 6922
rect 20328 5934 20374 5946
rect 20416 6320 20428 6330
rect 20462 6330 20468 6922
rect 20510 6928 20568 6934
rect 20510 6664 20522 6670
rect 20462 6320 20474 6330
rect 20416 5946 20428 5948
rect 20462 5946 20474 5948
rect 20416 5934 20474 5946
rect 20516 5946 20522 6664
rect 20556 6664 20568 6670
rect 20556 5946 20562 6664
rect 20596 6640 20630 6934
rect 20658 6928 20716 6934
rect 20658 6664 20670 6670
rect 20516 5934 20562 5946
rect 20590 6634 20636 6640
rect 20590 5946 20596 6634
rect 20630 5946 20636 6634
rect 20590 5812 20636 5946
rect 20664 5946 20670 6664
rect 20704 6664 20716 6670
rect 20758 6922 20804 6934
rect 20704 5946 20710 6664
rect 20758 6330 20764 6922
rect 20664 5934 20710 5946
rect 20752 6320 20764 6330
rect 20798 6330 20804 6922
rect 20846 6928 20904 6934
rect 20846 6664 20858 6670
rect 20798 6320 20810 6330
rect 20752 5946 20764 5948
rect 20798 5946 20810 5948
rect 20752 5934 20810 5946
rect 20852 5946 20858 6664
rect 20892 6664 20904 6670
rect 20892 5946 20898 6664
rect 20932 6640 20966 6934
rect 20994 6928 21052 6934
rect 20994 6664 21006 6670
rect 20852 5934 20898 5946
rect 20926 6634 20972 6640
rect 20926 5946 20932 6634
rect 20966 5946 20972 6634
rect 20926 5812 20972 5946
rect 21000 5946 21006 6664
rect 21040 6664 21052 6670
rect 21094 6922 21140 6934
rect 21040 5946 21046 6664
rect 21094 6330 21100 6922
rect 21000 5934 21046 5946
rect 21088 6320 21100 6330
rect 21134 6330 21140 6922
rect 21182 6928 21240 6934
rect 21182 6664 21194 6670
rect 21134 6320 21146 6330
rect 21088 5946 21100 5948
rect 21134 5946 21146 5948
rect 21088 5934 21146 5946
rect 21188 5946 21194 6664
rect 21228 6664 21240 6670
rect 21228 5946 21234 6664
rect 21268 6640 21302 6934
rect 21330 6928 21388 6934
rect 21330 6664 21342 6670
rect 21188 5934 21234 5946
rect 21262 6634 21308 6640
rect 21262 5946 21268 6634
rect 21302 5946 21308 6634
rect 21262 5812 21308 5946
rect 21336 5946 21342 6664
rect 21376 6664 21388 6670
rect 21430 6922 21476 6934
rect 21376 5946 21382 6664
rect 21430 6330 21436 6922
rect 21336 5934 21382 5946
rect 21424 6320 21436 6330
rect 21470 6330 21476 6922
rect 21518 6928 21576 6934
rect 21518 6664 21530 6670
rect 21470 6320 21482 6330
rect 21424 5946 21436 5948
rect 21470 5946 21482 5948
rect 21424 5934 21482 5946
rect 21524 5946 21530 6664
rect 21564 6664 21576 6670
rect 21564 5946 21570 6664
rect 21604 6640 21638 6934
rect 21666 6928 21724 6934
rect 21666 6664 21678 6670
rect 21524 5934 21570 5946
rect 21598 6634 21644 6640
rect 21598 5946 21604 6634
rect 21638 5946 21644 6634
rect 21598 5812 21644 5946
rect 21672 5946 21678 6664
rect 21712 6664 21724 6670
rect 21766 6922 21812 6934
rect 21712 5946 21718 6664
rect 21766 6330 21772 6922
rect 21672 5934 21718 5946
rect 21760 6320 21772 6330
rect 21806 6330 21812 6922
rect 21854 6928 21912 6934
rect 21854 6664 21866 6670
rect 21806 6320 21818 6330
rect 21760 5946 21772 5948
rect 21806 5946 21818 5948
rect 21760 5934 21818 5946
rect 21860 5946 21866 6664
rect 21900 6664 21912 6670
rect 21900 5946 21906 6664
rect 21940 6640 21996 6934
rect 21860 5934 21906 5946
rect 21934 6634 21996 6640
rect 21934 5946 21940 6634
rect 21974 5946 21996 6634
rect 21934 5812 21996 5946
rect 17426 5754 17454 5806
rect 17902 5754 17930 5806
rect 17426 5724 17930 5754
rect 19886 5806 22010 5812
rect 19886 5754 19906 5806
rect 21990 5754 22010 5806
rect 19886 5748 22010 5754
rect 15720 5494 15748 5662
rect 15804 5494 15832 5662
rect 15720 5484 15832 5494
rect 22090 5662 22202 7210
rect 28818 7122 28930 8704
rect 28958 8602 31454 8608
rect 28958 8550 28978 8602
rect 31434 8550 31454 8602
rect 28958 8544 31454 8550
rect 28958 8410 29070 8544
rect 29342 8410 29454 8544
rect 29746 8410 29858 8544
rect 30150 8410 30262 8544
rect 30554 8410 30666 8544
rect 30958 8410 31070 8544
rect 31342 8410 31454 8544
rect 28958 8398 29092 8410
rect 29174 8408 29220 8410
rect 28958 7422 28978 8398
rect 29012 7422 29052 8398
rect 29086 7422 29092 8398
rect 28958 7410 29092 7422
rect 29168 8398 29226 8408
rect 29168 7416 29226 7422
rect 29302 8398 29496 8410
rect 29578 8408 29624 8410
rect 29302 7422 29308 8398
rect 29342 7422 29382 8398
rect 29416 7422 29456 8398
rect 29490 7422 29496 8398
rect 29174 7410 29220 7416
rect 29302 7410 29496 7422
rect 29572 8398 29630 8408
rect 29572 7416 29630 7422
rect 29706 8398 29900 8410
rect 29982 8408 30028 8410
rect 29706 7422 29712 8398
rect 29746 7422 29786 8398
rect 29820 7422 29860 8398
rect 29894 7422 29900 8398
rect 29578 7410 29624 7416
rect 29706 7410 29900 7422
rect 29976 8398 30034 8408
rect 29976 7416 30034 7422
rect 30110 8398 30304 8410
rect 30386 8408 30432 8410
rect 30110 7422 30116 8398
rect 30150 7422 30190 8398
rect 30224 7422 30264 8398
rect 30298 7422 30304 8398
rect 29982 7410 30028 7416
rect 30110 7410 30304 7422
rect 30380 8398 30438 8408
rect 30380 7416 30438 7422
rect 30514 8398 30708 8410
rect 30790 8408 30836 8410
rect 30514 7422 30520 8398
rect 30554 7422 30594 8398
rect 30628 7422 30668 8398
rect 30702 7422 30708 8398
rect 30386 7410 30432 7416
rect 30514 7410 30708 7422
rect 30784 8398 30842 8408
rect 30784 7416 30842 7422
rect 30918 8398 31112 8410
rect 31194 8408 31240 8410
rect 30918 7422 30924 8398
rect 30958 7422 30998 8398
rect 31032 7422 31072 8398
rect 31106 7422 31112 8398
rect 30790 7410 30836 7416
rect 30918 7410 31112 7422
rect 31188 8398 31246 8408
rect 31188 7416 31246 7422
rect 31322 8398 31454 8410
rect 31322 7422 31328 8398
rect 31362 7422 31402 8398
rect 31436 7422 31454 8398
rect 31194 7410 31240 7416
rect 31322 7410 31454 7422
rect 29100 7363 29294 7370
rect 29100 7329 29114 7363
rect 29152 7329 29242 7363
rect 29280 7329 29294 7363
rect 29100 7310 29294 7329
rect 29504 7363 29698 7370
rect 29504 7329 29518 7363
rect 29556 7329 29646 7363
rect 29684 7329 29698 7363
rect 29504 7310 29698 7329
rect 29908 7363 30102 7370
rect 29908 7329 29922 7363
rect 29960 7329 30050 7363
rect 30088 7329 30102 7363
rect 29172 7268 29294 7310
rect 29172 7262 29422 7268
rect 29396 7210 29422 7262
rect 29172 7204 29422 7210
rect 28818 7064 28930 7070
rect 29288 7022 29422 7204
rect 29534 7128 29668 7310
rect 29908 7268 30102 7329
rect 30312 7363 30506 7370
rect 30312 7329 30326 7363
rect 30364 7329 30454 7363
rect 30492 7329 30506 7363
rect 29908 7262 30132 7268
rect 29908 7204 30132 7210
rect 29534 7122 29782 7128
rect 29758 7070 29782 7122
rect 29534 7064 29782 7070
rect 29288 7006 29446 7022
rect 29288 6972 29303 7006
rect 29337 6972 29397 7006
rect 29431 6972 29446 7006
rect 29288 6966 29446 6972
rect 29624 7006 29782 7064
rect 29624 6972 29639 7006
rect 29673 6972 29733 7006
rect 29767 6972 29782 7006
rect 29624 6966 29782 6972
rect 29960 7006 30118 7204
rect 30312 7128 30506 7329
rect 30716 7363 30910 7370
rect 30716 7329 30730 7363
rect 30768 7329 30858 7363
rect 30896 7329 30910 7363
rect 30716 7268 30910 7329
rect 30662 7262 30910 7268
rect 30886 7210 30910 7262
rect 30662 7204 30910 7210
rect 31120 7363 31314 7370
rect 31120 7329 31134 7363
rect 31172 7329 31262 7363
rect 31300 7329 31314 7363
rect 31120 7292 31314 7329
rect 30288 7122 30512 7128
rect 30288 7064 30512 7070
rect 29960 6972 29975 7006
rect 30009 6972 30069 7006
rect 30103 6972 30118 7006
rect 29960 6966 30118 6972
rect 30296 7006 30454 7064
rect 30662 7022 30774 7204
rect 31120 7128 31240 7292
rect 31008 7122 31240 7128
rect 31232 7070 31240 7122
rect 31008 7064 31240 7070
rect 31348 7262 31460 7268
rect 31008 7022 31126 7064
rect 30296 6972 30311 7006
rect 30345 6972 30405 7006
rect 30439 6972 30454 7006
rect 30296 6966 30454 6972
rect 30632 7006 30790 7022
rect 30632 6972 30647 7006
rect 30681 6972 30741 7006
rect 30775 6972 30790 7006
rect 30632 6966 30790 6972
rect 30968 7006 31126 7022
rect 30968 6972 30983 7006
rect 31017 6972 31077 7006
rect 31111 6972 31126 7006
rect 30968 6966 31126 6972
rect 23766 6614 24270 6664
rect 23766 6324 24028 6614
rect 24252 6324 24270 6614
rect 23766 5806 24270 6324
rect 29160 6642 29216 6934
rect 29244 6928 29302 6934
rect 29244 6664 29256 6670
rect 29160 6634 29222 6642
rect 29160 5946 29182 6634
rect 29216 5946 29222 6634
rect 29160 5812 29222 5946
rect 29250 5946 29256 6664
rect 29290 6664 29302 6670
rect 29344 6922 29390 6934
rect 29290 5946 29296 6664
rect 29344 6330 29350 6922
rect 29250 5934 29296 5946
rect 29338 6320 29350 6330
rect 29384 6330 29390 6922
rect 29432 6928 29490 6934
rect 29432 6664 29444 6670
rect 29384 6320 29396 6330
rect 29338 5946 29350 5948
rect 29384 5946 29396 5948
rect 29338 5934 29396 5946
rect 29438 5946 29444 6664
rect 29478 6664 29490 6670
rect 29478 5946 29484 6664
rect 29518 6640 29552 6934
rect 29580 6928 29638 6934
rect 29580 6664 29592 6670
rect 29438 5934 29484 5946
rect 29512 6634 29558 6640
rect 29512 5946 29518 6634
rect 29552 5946 29558 6634
rect 29512 5812 29558 5946
rect 29586 5946 29592 6664
rect 29626 6664 29638 6670
rect 29680 6922 29726 6934
rect 29626 5946 29632 6664
rect 29680 6330 29686 6922
rect 29586 5934 29632 5946
rect 29674 6320 29686 6330
rect 29720 6330 29726 6922
rect 29768 6928 29826 6934
rect 29768 6664 29780 6670
rect 29720 6320 29732 6330
rect 29674 5946 29686 5948
rect 29720 5946 29732 5948
rect 29674 5934 29732 5946
rect 29774 5946 29780 6664
rect 29814 6664 29826 6670
rect 29814 5946 29820 6664
rect 29854 6640 29888 6934
rect 29916 6928 29974 6934
rect 29916 6664 29928 6670
rect 29774 5934 29820 5946
rect 29848 6634 29894 6640
rect 29848 5946 29854 6634
rect 29888 5946 29894 6634
rect 29848 5812 29894 5946
rect 29922 5946 29928 6664
rect 29962 6664 29974 6670
rect 30016 6922 30062 6934
rect 29962 5946 29968 6664
rect 30016 6330 30022 6922
rect 29922 5934 29968 5946
rect 30010 6320 30022 6330
rect 30056 6330 30062 6922
rect 30104 6928 30162 6934
rect 30104 6664 30116 6670
rect 30056 6320 30068 6330
rect 30010 5946 30022 5948
rect 30056 5946 30068 5948
rect 30010 5934 30068 5946
rect 30110 5946 30116 6664
rect 30150 6664 30162 6670
rect 30150 5946 30156 6664
rect 30190 6640 30224 6934
rect 30252 6928 30310 6934
rect 30252 6664 30264 6670
rect 30110 5934 30156 5946
rect 30184 6634 30230 6640
rect 30184 5946 30190 6634
rect 30224 5946 30230 6634
rect 30184 5812 30230 5946
rect 30258 5946 30264 6664
rect 30298 6664 30310 6670
rect 30352 6922 30398 6934
rect 30298 5946 30304 6664
rect 30352 6330 30358 6922
rect 30258 5934 30304 5946
rect 30346 6320 30358 6330
rect 30392 6330 30398 6922
rect 30440 6928 30498 6934
rect 30440 6664 30452 6670
rect 30392 6320 30404 6330
rect 30346 5946 30358 5948
rect 30392 5946 30404 5948
rect 30346 5934 30404 5946
rect 30446 5946 30452 6664
rect 30486 6664 30498 6670
rect 30486 5946 30492 6664
rect 30526 6640 30560 6934
rect 30588 6928 30646 6934
rect 30588 6664 30600 6670
rect 30446 5934 30492 5946
rect 30520 6634 30566 6640
rect 30520 5946 30526 6634
rect 30560 5946 30566 6634
rect 30520 5812 30566 5946
rect 30594 5946 30600 6664
rect 30634 6664 30646 6670
rect 30688 6922 30734 6934
rect 30634 5946 30640 6664
rect 30688 6330 30694 6922
rect 30594 5934 30640 5946
rect 30682 6320 30694 6330
rect 30728 6330 30734 6922
rect 30776 6928 30834 6934
rect 30776 6664 30788 6670
rect 30728 6320 30740 6330
rect 30682 5946 30694 5948
rect 30728 5946 30740 5948
rect 30682 5934 30740 5946
rect 30782 5946 30788 6664
rect 30822 6664 30834 6670
rect 30822 5946 30828 6664
rect 30862 6640 30896 6934
rect 30924 6928 30982 6934
rect 30924 6664 30936 6670
rect 30782 5934 30828 5946
rect 30856 6634 30902 6640
rect 30856 5946 30862 6634
rect 30896 5946 30902 6634
rect 30856 5812 30902 5946
rect 30930 5946 30936 6664
rect 30970 6664 30982 6670
rect 31024 6922 31070 6934
rect 30970 5946 30976 6664
rect 31024 6330 31030 6922
rect 30930 5934 30976 5946
rect 31018 6320 31030 6330
rect 31064 6330 31070 6922
rect 31112 6928 31170 6934
rect 31112 6664 31124 6670
rect 31064 6320 31076 6330
rect 31018 5946 31030 5948
rect 31064 5946 31076 5948
rect 31018 5934 31076 5946
rect 31118 5946 31124 6664
rect 31158 6664 31170 6670
rect 31158 5946 31164 6664
rect 31198 6640 31254 6934
rect 31118 5934 31164 5946
rect 31192 6634 31254 6640
rect 31192 5946 31198 6634
rect 31232 5946 31254 6634
rect 31192 5812 31254 5946
rect 23766 5754 23794 5806
rect 24242 5754 24270 5806
rect 23766 5724 24270 5754
rect 29144 5806 31268 5812
rect 29144 5754 29164 5806
rect 31248 5754 31268 5806
rect 29144 5748 31268 5754
rect 22090 5494 22118 5662
rect 22174 5494 22202 5662
rect 22090 5484 22202 5494
rect 31348 5662 31460 7210
rect 31348 5494 31376 5662
rect 31432 5494 31460 5662
rect 31348 5484 31460 5494
rect -2418 5434 -2306 5444
<< via1 >>
rect -4918 8654 -4862 8822
rect 480 8704 536 8872
rect -4788 8500 -2312 8552
rect -4598 7372 -4586 8348
rect -4586 7372 -4552 8348
rect -4552 7372 -4540 8348
rect -4194 7372 -4182 8348
rect -4182 7372 -4148 8348
rect -4148 7372 -4136 8348
rect -3790 7372 -3778 8348
rect -3778 7372 -3744 8348
rect -3744 7372 -3732 8348
rect -3386 7372 -3374 8348
rect -3374 7372 -3340 8348
rect -3340 7372 -3328 8348
rect -2982 7372 -2970 8348
rect -2970 7372 -2936 8348
rect -2936 7372 -2924 8348
rect -2578 7372 -2566 8348
rect -2566 7372 -2532 8348
rect -2532 7372 -2520 8348
rect -4594 7160 -4370 7212
rect -4948 7020 -4836 7072
rect -3858 7160 -3634 7212
rect -4232 7020 -4008 7072
rect -3104 7160 -2880 7212
rect -3478 7020 -3254 7072
rect -2758 7020 -2534 7072
rect -2418 7160 -2306 7212
rect -5226 6326 -5002 6616
rect -4428 6872 -4370 6874
rect -4428 5898 -4416 6872
rect -4416 5898 -4382 6872
rect -4382 5898 -4370 6872
rect -4092 6872 -4034 6874
rect -4092 5898 -4080 6872
rect -4080 5898 -4046 6872
rect -4046 5898 -4034 6872
rect -3756 6872 -3698 6874
rect -3756 5898 -3744 6872
rect -3744 5898 -3710 6872
rect -3710 5898 -3698 6872
rect -3420 6872 -3362 6874
rect -3420 5898 -3408 6872
rect -3408 5898 -3374 6872
rect -3374 5898 -3362 6872
rect -3084 6872 -3026 6874
rect -3084 5898 -3072 6872
rect -3072 5898 -3038 6872
rect -3038 5898 -3026 6872
rect -2748 6872 -2690 6874
rect -2748 5898 -2736 6872
rect -2736 5898 -2702 6872
rect -2702 5898 -2690 6872
rect -5200 5704 -2518 5756
rect 6850 8704 6906 8872
rect 610 8550 3066 8602
rect 800 7422 812 8398
rect 812 7422 846 8398
rect 846 7422 858 8398
rect 1204 7422 1216 8398
rect 1216 7422 1250 8398
rect 1250 7422 1262 8398
rect 1608 7422 1620 8398
rect 1620 7422 1654 8398
rect 1654 7422 1666 8398
rect 2012 7422 2024 8398
rect 2024 7422 2058 8398
rect 2058 7422 2070 8398
rect 2416 7422 2428 8398
rect 2428 7422 2462 8398
rect 2462 7422 2474 8398
rect 2820 7422 2832 8398
rect 2832 7422 2866 8398
rect 2866 7422 2878 8398
rect 804 7210 1028 7262
rect 450 7070 562 7122
rect 1540 7210 1764 7262
rect 1166 7070 1390 7122
rect 2294 7210 2518 7262
rect 1920 7070 2144 7122
rect 2640 7070 2864 7122
rect 2980 7210 3092 7262
rect -1422 6324 -1198 6614
rect 876 6922 934 6928
rect 876 6670 888 6922
rect 888 6670 922 6922
rect 922 6670 934 6922
rect 1064 6922 1122 6928
rect 1064 6670 1076 6922
rect 1076 6670 1110 6922
rect 1110 6670 1122 6922
rect 970 5948 982 6320
rect 982 5948 1016 6320
rect 1016 5948 1028 6320
rect 1212 6922 1270 6928
rect 1212 6670 1224 6922
rect 1224 6670 1258 6922
rect 1258 6670 1270 6922
rect 1400 6922 1458 6928
rect 1400 6670 1412 6922
rect 1412 6670 1446 6922
rect 1446 6670 1458 6922
rect 1306 5948 1318 6320
rect 1318 5948 1352 6320
rect 1352 5948 1364 6320
rect 1548 6922 1606 6928
rect 1548 6670 1560 6922
rect 1560 6670 1594 6922
rect 1594 6670 1606 6922
rect 1736 6922 1794 6928
rect 1736 6670 1748 6922
rect 1748 6670 1782 6922
rect 1782 6670 1794 6922
rect 1642 5948 1654 6320
rect 1654 5948 1688 6320
rect 1688 5948 1700 6320
rect 1884 6922 1942 6928
rect 1884 6670 1896 6922
rect 1896 6670 1930 6922
rect 1930 6670 1942 6922
rect 2072 6922 2130 6928
rect 2072 6670 2084 6922
rect 2084 6670 2118 6922
rect 2118 6670 2130 6922
rect 1978 5948 1990 6320
rect 1990 5948 2024 6320
rect 2024 5948 2036 6320
rect 2220 6922 2278 6928
rect 2220 6670 2232 6922
rect 2232 6670 2266 6922
rect 2266 6670 2278 6922
rect 2408 6922 2466 6928
rect 2408 6670 2420 6922
rect 2420 6670 2454 6922
rect 2454 6670 2466 6922
rect 2314 5948 2326 6320
rect 2326 5948 2360 6320
rect 2360 5948 2372 6320
rect 2556 6922 2614 6928
rect 2556 6670 2568 6922
rect 2568 6670 2602 6922
rect 2602 6670 2614 6922
rect 2744 6922 2802 6928
rect 2744 6670 2756 6922
rect 2756 6670 2790 6922
rect 2790 6670 2802 6922
rect 2650 5948 2662 6320
rect 2662 5948 2696 6320
rect 2696 5948 2708 6320
rect -1656 5754 -1208 5806
rect 796 5754 2880 5806
rect -2390 5444 -2334 5612
rect 13220 8704 13276 8872
rect 6980 8550 9436 8602
rect 7170 7422 7182 8398
rect 7182 7422 7216 8398
rect 7216 7422 7228 8398
rect 7574 7422 7586 8398
rect 7586 7422 7620 8398
rect 7620 7422 7632 8398
rect 7978 7422 7990 8398
rect 7990 7422 8024 8398
rect 8024 7422 8036 8398
rect 8382 7422 8394 8398
rect 8394 7422 8428 8398
rect 8428 7422 8440 8398
rect 8786 7422 8798 8398
rect 8798 7422 8832 8398
rect 8832 7422 8844 8398
rect 9190 7422 9202 8398
rect 9202 7422 9236 8398
rect 9236 7422 9248 8398
rect 7174 7210 7398 7262
rect 6820 7070 6932 7122
rect 7910 7210 8134 7262
rect 7536 7070 7760 7122
rect 8664 7210 8888 7262
rect 8290 7070 8514 7122
rect 9010 7070 9234 7122
rect 9350 7210 9462 7262
rect 4948 6324 5172 6614
rect 7246 6922 7304 6928
rect 7246 6670 7258 6922
rect 7258 6670 7292 6922
rect 7292 6670 7304 6922
rect 7434 6922 7492 6928
rect 7434 6670 7446 6922
rect 7446 6670 7480 6922
rect 7480 6670 7492 6922
rect 7340 5948 7352 6320
rect 7352 5948 7386 6320
rect 7386 5948 7398 6320
rect 7582 6922 7640 6928
rect 7582 6670 7594 6922
rect 7594 6670 7628 6922
rect 7628 6670 7640 6922
rect 7770 6922 7828 6928
rect 7770 6670 7782 6922
rect 7782 6670 7816 6922
rect 7816 6670 7828 6922
rect 7676 5948 7688 6320
rect 7688 5948 7722 6320
rect 7722 5948 7734 6320
rect 7918 6922 7976 6928
rect 7918 6670 7930 6922
rect 7930 6670 7964 6922
rect 7964 6670 7976 6922
rect 8106 6922 8164 6928
rect 8106 6670 8118 6922
rect 8118 6670 8152 6922
rect 8152 6670 8164 6922
rect 8012 5948 8024 6320
rect 8024 5948 8058 6320
rect 8058 5948 8070 6320
rect 8254 6922 8312 6928
rect 8254 6670 8266 6922
rect 8266 6670 8300 6922
rect 8300 6670 8312 6922
rect 8442 6922 8500 6928
rect 8442 6670 8454 6922
rect 8454 6670 8488 6922
rect 8488 6670 8500 6922
rect 8348 5948 8360 6320
rect 8360 5948 8394 6320
rect 8394 5948 8406 6320
rect 8590 6922 8648 6928
rect 8590 6670 8602 6922
rect 8602 6670 8636 6922
rect 8636 6670 8648 6922
rect 8778 6922 8836 6928
rect 8778 6670 8790 6922
rect 8790 6670 8824 6922
rect 8824 6670 8836 6922
rect 8684 5948 8696 6320
rect 8696 5948 8730 6320
rect 8730 5948 8742 6320
rect 8926 6922 8984 6928
rect 8926 6670 8938 6922
rect 8938 6670 8972 6922
rect 8972 6670 8984 6922
rect 9114 6922 9172 6928
rect 9114 6670 9126 6922
rect 9126 6670 9160 6922
rect 9160 6670 9172 6922
rect 9020 5948 9032 6320
rect 9032 5948 9066 6320
rect 9066 5948 9078 6320
rect 4714 5754 5162 5806
rect 7166 5754 9250 5806
rect 3008 5494 3064 5662
rect 19590 8704 19646 8872
rect 13350 8550 15806 8602
rect 13540 7422 13552 8398
rect 13552 7422 13586 8398
rect 13586 7422 13598 8398
rect 13944 7422 13956 8398
rect 13956 7422 13990 8398
rect 13990 7422 14002 8398
rect 14348 7422 14360 8398
rect 14360 7422 14394 8398
rect 14394 7422 14406 8398
rect 14752 7422 14764 8398
rect 14764 7422 14798 8398
rect 14798 7422 14810 8398
rect 15156 7422 15168 8398
rect 15168 7422 15202 8398
rect 15202 7422 15214 8398
rect 15560 7422 15572 8398
rect 15572 7422 15606 8398
rect 15606 7422 15618 8398
rect 13544 7210 13768 7262
rect 13190 7070 13302 7122
rect 14280 7210 14504 7262
rect 13906 7070 14130 7122
rect 15034 7210 15258 7262
rect 14660 7070 14884 7122
rect 15380 7070 15604 7122
rect 15720 7210 15832 7262
rect 11318 6324 11542 6614
rect 13616 6922 13674 6928
rect 13616 6670 13628 6922
rect 13628 6670 13662 6922
rect 13662 6670 13674 6922
rect 13804 6922 13862 6928
rect 13804 6670 13816 6922
rect 13816 6670 13850 6922
rect 13850 6670 13862 6922
rect 13710 5948 13722 6320
rect 13722 5948 13756 6320
rect 13756 5948 13768 6320
rect 13952 6922 14010 6928
rect 13952 6670 13964 6922
rect 13964 6670 13998 6922
rect 13998 6670 14010 6922
rect 14140 6922 14198 6928
rect 14140 6670 14152 6922
rect 14152 6670 14186 6922
rect 14186 6670 14198 6922
rect 14046 5948 14058 6320
rect 14058 5948 14092 6320
rect 14092 5948 14104 6320
rect 14288 6922 14346 6928
rect 14288 6670 14300 6922
rect 14300 6670 14334 6922
rect 14334 6670 14346 6922
rect 14476 6922 14534 6928
rect 14476 6670 14488 6922
rect 14488 6670 14522 6922
rect 14522 6670 14534 6922
rect 14382 5948 14394 6320
rect 14394 5948 14428 6320
rect 14428 5948 14440 6320
rect 14624 6922 14682 6928
rect 14624 6670 14636 6922
rect 14636 6670 14670 6922
rect 14670 6670 14682 6922
rect 14812 6922 14870 6928
rect 14812 6670 14824 6922
rect 14824 6670 14858 6922
rect 14858 6670 14870 6922
rect 14718 5948 14730 6320
rect 14730 5948 14764 6320
rect 14764 5948 14776 6320
rect 14960 6922 15018 6928
rect 14960 6670 14972 6922
rect 14972 6670 15006 6922
rect 15006 6670 15018 6922
rect 15148 6922 15206 6928
rect 15148 6670 15160 6922
rect 15160 6670 15194 6922
rect 15194 6670 15206 6922
rect 15054 5948 15066 6320
rect 15066 5948 15100 6320
rect 15100 5948 15112 6320
rect 15296 6922 15354 6928
rect 15296 6670 15308 6922
rect 15308 6670 15342 6922
rect 15342 6670 15354 6922
rect 15484 6922 15542 6928
rect 15484 6670 15496 6922
rect 15496 6670 15530 6922
rect 15530 6670 15542 6922
rect 15390 5948 15402 6320
rect 15402 5948 15436 6320
rect 15436 5948 15448 6320
rect 11084 5754 11532 5806
rect 13536 5754 15620 5806
rect 9378 5494 9434 5662
rect 28848 8704 28904 8872
rect 19720 8550 22176 8602
rect 19910 7422 19922 8398
rect 19922 7422 19956 8398
rect 19956 7422 19968 8398
rect 20314 7422 20326 8398
rect 20326 7422 20360 8398
rect 20360 7422 20372 8398
rect 20718 7422 20730 8398
rect 20730 7422 20764 8398
rect 20764 7422 20776 8398
rect 21122 7422 21134 8398
rect 21134 7422 21168 8398
rect 21168 7422 21180 8398
rect 21526 7422 21538 8398
rect 21538 7422 21572 8398
rect 21572 7422 21584 8398
rect 21930 7422 21942 8398
rect 21942 7422 21976 8398
rect 21976 7422 21988 8398
rect 19914 7210 20138 7262
rect 19560 7070 19672 7122
rect 20650 7210 20874 7262
rect 20276 7070 20500 7122
rect 21404 7210 21628 7262
rect 21030 7070 21254 7122
rect 21750 7070 21974 7122
rect 22090 7210 22202 7262
rect 17688 6324 17912 6614
rect 19986 6922 20044 6928
rect 19986 6670 19998 6922
rect 19998 6670 20032 6922
rect 20032 6670 20044 6922
rect 20174 6922 20232 6928
rect 20174 6670 20186 6922
rect 20186 6670 20220 6922
rect 20220 6670 20232 6922
rect 20080 5948 20092 6320
rect 20092 5948 20126 6320
rect 20126 5948 20138 6320
rect 20322 6922 20380 6928
rect 20322 6670 20334 6922
rect 20334 6670 20368 6922
rect 20368 6670 20380 6922
rect 20510 6922 20568 6928
rect 20510 6670 20522 6922
rect 20522 6670 20556 6922
rect 20556 6670 20568 6922
rect 20416 5948 20428 6320
rect 20428 5948 20462 6320
rect 20462 5948 20474 6320
rect 20658 6922 20716 6928
rect 20658 6670 20670 6922
rect 20670 6670 20704 6922
rect 20704 6670 20716 6922
rect 20846 6922 20904 6928
rect 20846 6670 20858 6922
rect 20858 6670 20892 6922
rect 20892 6670 20904 6922
rect 20752 5948 20764 6320
rect 20764 5948 20798 6320
rect 20798 5948 20810 6320
rect 20994 6922 21052 6928
rect 20994 6670 21006 6922
rect 21006 6670 21040 6922
rect 21040 6670 21052 6922
rect 21182 6922 21240 6928
rect 21182 6670 21194 6922
rect 21194 6670 21228 6922
rect 21228 6670 21240 6922
rect 21088 5948 21100 6320
rect 21100 5948 21134 6320
rect 21134 5948 21146 6320
rect 21330 6922 21388 6928
rect 21330 6670 21342 6922
rect 21342 6670 21376 6922
rect 21376 6670 21388 6922
rect 21518 6922 21576 6928
rect 21518 6670 21530 6922
rect 21530 6670 21564 6922
rect 21564 6670 21576 6922
rect 21424 5948 21436 6320
rect 21436 5948 21470 6320
rect 21470 5948 21482 6320
rect 21666 6922 21724 6928
rect 21666 6670 21678 6922
rect 21678 6670 21712 6922
rect 21712 6670 21724 6922
rect 21854 6922 21912 6928
rect 21854 6670 21866 6922
rect 21866 6670 21900 6922
rect 21900 6670 21912 6922
rect 21760 5948 21772 6320
rect 21772 5948 21806 6320
rect 21806 5948 21818 6320
rect 17454 5754 17902 5806
rect 19906 5754 21990 5806
rect 15748 5494 15804 5662
rect 28978 8550 31434 8602
rect 29168 7422 29180 8398
rect 29180 7422 29214 8398
rect 29214 7422 29226 8398
rect 29572 7422 29584 8398
rect 29584 7422 29618 8398
rect 29618 7422 29630 8398
rect 29976 7422 29988 8398
rect 29988 7422 30022 8398
rect 30022 7422 30034 8398
rect 30380 7422 30392 8398
rect 30392 7422 30426 8398
rect 30426 7422 30438 8398
rect 30784 7422 30796 8398
rect 30796 7422 30830 8398
rect 30830 7422 30842 8398
rect 31188 7422 31200 8398
rect 31200 7422 31234 8398
rect 31234 7422 31246 8398
rect 29172 7210 29396 7262
rect 28818 7070 28930 7122
rect 29908 7210 30132 7262
rect 29534 7070 29758 7122
rect 30662 7210 30886 7262
rect 30288 7070 30512 7122
rect 31008 7070 31232 7122
rect 31348 7210 31460 7262
rect 24028 6324 24252 6614
rect 29244 6922 29302 6928
rect 29244 6670 29256 6922
rect 29256 6670 29290 6922
rect 29290 6670 29302 6922
rect 29432 6922 29490 6928
rect 29432 6670 29444 6922
rect 29444 6670 29478 6922
rect 29478 6670 29490 6922
rect 29338 5948 29350 6320
rect 29350 5948 29384 6320
rect 29384 5948 29396 6320
rect 29580 6922 29638 6928
rect 29580 6670 29592 6922
rect 29592 6670 29626 6922
rect 29626 6670 29638 6922
rect 29768 6922 29826 6928
rect 29768 6670 29780 6922
rect 29780 6670 29814 6922
rect 29814 6670 29826 6922
rect 29674 5948 29686 6320
rect 29686 5948 29720 6320
rect 29720 5948 29732 6320
rect 29916 6922 29974 6928
rect 29916 6670 29928 6922
rect 29928 6670 29962 6922
rect 29962 6670 29974 6922
rect 30104 6922 30162 6928
rect 30104 6670 30116 6922
rect 30116 6670 30150 6922
rect 30150 6670 30162 6922
rect 30010 5948 30022 6320
rect 30022 5948 30056 6320
rect 30056 5948 30068 6320
rect 30252 6922 30310 6928
rect 30252 6670 30264 6922
rect 30264 6670 30298 6922
rect 30298 6670 30310 6922
rect 30440 6922 30498 6928
rect 30440 6670 30452 6922
rect 30452 6670 30486 6922
rect 30486 6670 30498 6922
rect 30346 5948 30358 6320
rect 30358 5948 30392 6320
rect 30392 5948 30404 6320
rect 30588 6922 30646 6928
rect 30588 6670 30600 6922
rect 30600 6670 30634 6922
rect 30634 6670 30646 6922
rect 30776 6922 30834 6928
rect 30776 6670 30788 6922
rect 30788 6670 30822 6922
rect 30822 6670 30834 6922
rect 30682 5948 30694 6320
rect 30694 5948 30728 6320
rect 30728 5948 30740 6320
rect 30924 6922 30982 6928
rect 30924 6670 30936 6922
rect 30936 6670 30970 6922
rect 30970 6670 30982 6922
rect 31112 6922 31170 6928
rect 31112 6670 31124 6922
rect 31124 6670 31158 6922
rect 31158 6670 31170 6922
rect 31018 5948 31030 6320
rect 31030 5948 31064 6320
rect 31064 5948 31076 6320
rect 23794 5754 24242 5806
rect 29164 5754 31248 5806
rect 22118 5494 22174 5662
rect 31376 5494 31432 5662
<< metal2 >>
rect 450 8872 562 8882
rect -4948 8822 -4836 8832
rect -4948 8654 -4918 8822
rect -4862 8654 -4836 8822
rect 450 8704 480 8872
rect 536 8704 562 8872
rect 6820 8872 6932 8882
rect 450 8694 562 8704
rect -4948 8644 -4836 8654
rect -4808 8580 -1982 8694
rect -4808 8552 -2212 8580
rect -4808 8500 -4788 8552
rect -2312 8500 -2212 8552
rect -4808 8414 -2212 8500
rect -4598 8348 -4540 8358
rect -4598 7360 -4540 7372
rect -4194 8348 -4136 8358
rect -4194 7360 -4136 7372
rect -3790 8348 -3732 8358
rect -3790 7360 -3732 7372
rect -3386 8348 -3328 8358
rect -3386 7360 -3328 7372
rect -2982 8348 -2924 8358
rect -2982 7360 -2924 7372
rect -2578 8348 -2520 8358
rect -2578 7360 -2520 7372
rect -4594 7242 -4472 7270
rect -4672 7212 -2306 7242
rect -4672 7160 -4594 7212
rect -4370 7160 -3858 7212
rect -3634 7160 -3104 7212
rect -2880 7160 -2418 7212
rect -4672 7130 -2306 7160
rect -4948 7072 -2446 7102
rect -4836 7020 -4232 7072
rect -4008 7020 -3478 7072
rect -3254 7020 -2758 7072
rect -2534 7020 -2446 7072
rect -4948 6990 -2446 7020
rect -4428 6874 -4370 6886
rect -5242 6616 -4984 6632
rect -5242 6326 -5226 6616
rect -5002 6326 -4984 6616
rect -5242 6306 -4984 6326
rect -4428 5884 -4370 5898
rect -4092 6874 -4034 6886
rect -4092 5884 -4034 5898
rect -3756 6874 -3698 6886
rect -3756 5884 -3698 5898
rect -3420 6874 -3362 6886
rect -3420 5884 -3362 5898
rect -3084 6874 -3026 6886
rect -3084 5884 -3026 5898
rect -2748 6874 -2690 6886
rect -2224 6722 -2212 8414
rect -1994 6722 -1982 8580
rect 590 8602 3788 8716
rect 6820 8704 6850 8872
rect 6906 8704 6932 8872
rect 13190 8872 13302 8882
rect 6820 8694 6932 8704
rect 590 8550 610 8602
rect 3066 8580 3788 8602
rect 3066 8550 3572 8580
rect 590 8436 3572 8550
rect 800 8398 858 8408
rect 800 7410 858 7422
rect 1204 8398 1262 8408
rect 1204 7410 1262 7422
rect 1608 8398 1666 8408
rect 1608 7410 1666 7422
rect 2012 8398 2070 8408
rect 2012 7410 2070 7422
rect 2416 8398 2474 8408
rect 2416 7410 2474 7422
rect 2820 8398 2878 8408
rect 2820 7410 2878 7422
rect 804 7292 926 7320
rect 726 7262 3092 7292
rect 726 7210 804 7262
rect 1028 7210 1540 7262
rect 1764 7210 2294 7262
rect 2518 7210 2980 7262
rect 726 7180 3092 7210
rect 450 7122 2952 7152
rect 562 7070 1166 7122
rect 1390 7070 1920 7122
rect 2144 7070 2640 7122
rect 2864 7070 2952 7122
rect 450 7040 2952 7070
rect -2224 6710 -1982 6722
rect -1684 6928 2802 6934
rect -1684 6884 876 6928
rect -1684 6772 -1640 6884
rect -646 6772 876 6884
rect -1684 6710 876 6772
rect 934 6710 1064 6928
rect 876 6664 934 6670
rect 1122 6710 1212 6928
rect 1064 6664 1122 6670
rect 1270 6710 1400 6928
rect 1212 6664 1270 6670
rect 1458 6710 1548 6928
rect 1400 6664 1458 6670
rect 1606 6710 1736 6928
rect 1548 6664 1606 6670
rect 1794 6710 1884 6928
rect 1736 6664 1794 6670
rect 1942 6710 2072 6928
rect 1884 6664 1942 6670
rect 2130 6710 2220 6928
rect 2072 6664 2130 6670
rect 2278 6710 2408 6928
rect 2220 6664 2278 6670
rect 2466 6710 2556 6928
rect 2408 6664 2466 6670
rect 2614 6710 2744 6928
rect 2556 6664 2614 6670
rect 3516 6728 3572 8436
rect 3684 6728 3788 8580
rect 6960 8602 10158 8716
rect 13190 8704 13220 8872
rect 13276 8704 13302 8872
rect 19560 8872 19672 8882
rect 13190 8694 13302 8704
rect 6960 8550 6980 8602
rect 9436 8580 10158 8602
rect 9436 8550 9942 8580
rect 6960 8436 9942 8550
rect 7170 8398 7228 8408
rect 7170 7410 7228 7422
rect 7574 8398 7632 8408
rect 7574 7410 7632 7422
rect 7978 8398 8036 8408
rect 7978 7410 8036 7422
rect 8382 8398 8440 8408
rect 8382 7410 8440 7422
rect 8786 8398 8844 8408
rect 8786 7410 8844 7422
rect 9190 8398 9248 8408
rect 9190 7410 9248 7422
rect 7174 7292 7296 7320
rect 7096 7262 9462 7292
rect 7096 7210 7174 7262
rect 7398 7210 7910 7262
rect 8134 7210 8664 7262
rect 8888 7210 9350 7262
rect 7096 7180 9462 7210
rect 6820 7122 9322 7152
rect 6932 7070 7536 7122
rect 7760 7070 8290 7122
rect 8514 7070 9010 7122
rect 9234 7070 9322 7122
rect 6820 7040 9322 7070
rect 3516 6710 3788 6728
rect 4686 6928 9172 6934
rect 4686 6884 7246 6928
rect 4686 6772 4730 6884
rect 5724 6772 7246 6884
rect 4686 6710 7246 6772
rect 2744 6664 2802 6670
rect 7304 6710 7434 6928
rect 7246 6664 7304 6670
rect 7492 6710 7582 6928
rect 7434 6664 7492 6670
rect 7640 6710 7770 6928
rect 7582 6664 7640 6670
rect 7828 6710 7918 6928
rect 7770 6664 7828 6670
rect 7976 6710 8106 6928
rect 7918 6664 7976 6670
rect 8164 6710 8254 6928
rect 8106 6664 8164 6670
rect 8312 6710 8442 6928
rect 8254 6664 8312 6670
rect 8500 6710 8590 6928
rect 8442 6664 8500 6670
rect 8648 6710 8778 6928
rect 8590 6664 8648 6670
rect 8836 6710 8926 6928
rect 8778 6664 8836 6670
rect 8984 6710 9114 6928
rect 8926 6664 8984 6670
rect 9886 6728 9942 8436
rect 10054 6728 10158 8580
rect 13330 8602 16528 8716
rect 19560 8704 19590 8872
rect 19646 8704 19672 8872
rect 28818 8872 28930 8882
rect 19560 8694 19672 8704
rect 13330 8550 13350 8602
rect 15806 8580 16528 8602
rect 15806 8550 16312 8580
rect 13330 8436 16312 8550
rect 13540 8398 13598 8408
rect 13540 7410 13598 7422
rect 13944 8398 14002 8408
rect 13944 7410 14002 7422
rect 14348 8398 14406 8408
rect 14348 7410 14406 7422
rect 14752 8398 14810 8408
rect 14752 7410 14810 7422
rect 15156 8398 15214 8408
rect 15156 7410 15214 7422
rect 15560 8398 15618 8408
rect 15560 7410 15618 7422
rect 13544 7292 13666 7320
rect 13466 7262 15832 7292
rect 13466 7210 13544 7262
rect 13768 7210 14280 7262
rect 14504 7210 15034 7262
rect 15258 7210 15720 7262
rect 13466 7180 15832 7210
rect 13190 7122 15692 7152
rect 13302 7070 13906 7122
rect 14130 7070 14660 7122
rect 14884 7070 15380 7122
rect 15604 7070 15692 7122
rect 13190 7040 15692 7070
rect 9886 6710 10158 6728
rect 11056 6928 15542 6934
rect 11056 6884 13616 6928
rect 11056 6772 11100 6884
rect 12094 6772 13616 6884
rect 11056 6710 13616 6772
rect 9114 6664 9172 6670
rect 13674 6710 13804 6928
rect 13616 6664 13674 6670
rect 13862 6710 13952 6928
rect 13804 6664 13862 6670
rect 14010 6710 14140 6928
rect 13952 6664 14010 6670
rect 14198 6710 14288 6928
rect 14140 6664 14198 6670
rect 14346 6710 14476 6928
rect 14288 6664 14346 6670
rect 14534 6710 14624 6928
rect 14476 6664 14534 6670
rect 14682 6710 14812 6928
rect 14624 6664 14682 6670
rect 14870 6710 14960 6928
rect 14812 6664 14870 6670
rect 15018 6710 15148 6928
rect 14960 6664 15018 6670
rect 15206 6710 15296 6928
rect 15148 6664 15206 6670
rect 15354 6710 15484 6928
rect 15296 6664 15354 6670
rect 16256 6728 16312 8436
rect 16424 6728 16528 8580
rect 19700 8602 22898 8716
rect 28818 8704 28848 8872
rect 28904 8704 28930 8872
rect 28818 8694 28930 8704
rect 19700 8550 19720 8602
rect 22176 8580 22898 8602
rect 22176 8550 22682 8580
rect 19700 8436 22682 8550
rect 19910 8398 19968 8408
rect 19910 7410 19968 7422
rect 20314 8398 20372 8408
rect 20314 7410 20372 7422
rect 20718 8398 20776 8408
rect 20718 7410 20776 7422
rect 21122 8398 21180 8408
rect 21122 7410 21180 7422
rect 21526 8398 21584 8408
rect 21526 7410 21584 7422
rect 21930 8398 21988 8408
rect 21930 7410 21988 7422
rect 19914 7292 20036 7320
rect 19836 7262 22202 7292
rect 19836 7210 19914 7262
rect 20138 7210 20650 7262
rect 20874 7210 21404 7262
rect 21628 7210 22090 7262
rect 19836 7180 22202 7210
rect 19560 7122 22062 7152
rect 19672 7070 20276 7122
rect 20500 7070 21030 7122
rect 21254 7070 21750 7122
rect 21974 7070 22062 7122
rect 19560 7040 22062 7070
rect 16256 6710 16528 6728
rect 17426 6928 21912 6934
rect 17426 6884 19986 6928
rect 17426 6772 17470 6884
rect 18464 6772 19986 6884
rect 17426 6710 19986 6772
rect 15484 6664 15542 6670
rect 20044 6710 20174 6928
rect 19986 6664 20044 6670
rect 20232 6710 20322 6928
rect 20174 6664 20232 6670
rect 20380 6710 20510 6928
rect 20322 6664 20380 6670
rect 20568 6710 20658 6928
rect 20510 6664 20568 6670
rect 20716 6710 20846 6928
rect 20658 6664 20716 6670
rect 20904 6710 20994 6928
rect 20846 6664 20904 6670
rect 21052 6710 21182 6928
rect 20994 6664 21052 6670
rect 21240 6710 21330 6928
rect 21182 6664 21240 6670
rect 21388 6710 21518 6928
rect 21330 6664 21388 6670
rect 21576 6710 21666 6928
rect 21518 6664 21576 6670
rect 21724 6710 21854 6928
rect 21666 6664 21724 6670
rect 22626 6728 22682 8436
rect 22794 6728 22898 8580
rect 28958 8602 35980 8828
rect 28958 8550 28978 8602
rect 31434 8550 35980 8602
rect 28958 8480 35980 8550
rect 28958 8436 35668 8480
rect 29168 8398 29226 8408
rect 29168 7410 29226 7422
rect 29572 8398 29630 8408
rect 29572 7410 29630 7422
rect 29976 8398 30034 8408
rect 29976 7410 30034 7422
rect 30380 8398 30438 8408
rect 30380 7410 30438 7422
rect 30784 8398 30842 8408
rect 30784 7410 30842 7422
rect 31188 8398 31246 8408
rect 31188 7410 31246 7422
rect 29172 7292 29294 7320
rect 29094 7262 31460 7292
rect 29094 7210 29172 7262
rect 29396 7210 29908 7262
rect 30132 7210 30662 7262
rect 30886 7210 31348 7262
rect 29094 7180 31460 7210
rect 28818 7122 31320 7152
rect 28930 7070 29534 7122
rect 29758 7070 30288 7122
rect 30512 7070 31008 7122
rect 31232 7070 31320 7122
rect 28818 7040 31320 7070
rect 22626 6710 22898 6728
rect 23766 6928 31170 6934
rect 23766 6884 29244 6928
rect 23766 6772 23810 6884
rect 24804 6772 29244 6884
rect 23766 6710 29244 6772
rect 21854 6664 21912 6670
rect 29160 6670 29244 6710
rect 29302 6670 29432 6928
rect 29490 6670 29580 6928
rect 29638 6670 29768 6928
rect 29826 6670 29916 6928
rect 29974 6670 30104 6928
rect 30162 6670 30252 6928
rect 30310 6670 30440 6928
rect 30498 6670 30588 6928
rect 30646 6670 30776 6928
rect 30834 6670 30924 6928
rect 30982 6670 31112 6928
rect -1438 6614 -1180 6630
rect -1438 6324 -1422 6614
rect -1198 6324 -1180 6614
rect 4932 6614 5190 6630
rect -1438 6304 -1180 6324
rect 970 6320 1028 6330
rect 970 5934 1028 5948
rect 1306 6320 1364 6330
rect 1306 5934 1364 5948
rect 1642 6320 1700 6330
rect 1642 5934 1700 5948
rect 1978 6320 2036 6330
rect 1978 5934 2036 5948
rect 2314 6320 2372 6330
rect 2314 5934 2372 5948
rect 2650 6320 2708 6330
rect 4932 6324 4948 6614
rect 5172 6324 5190 6614
rect 11302 6614 11560 6630
rect 4932 6304 5190 6324
rect 7340 6320 7398 6330
rect 2650 5934 2708 5948
rect 7340 5934 7398 5948
rect 7676 6320 7734 6330
rect 7676 5934 7734 5948
rect 8012 6320 8070 6330
rect 8012 5934 8070 5948
rect 8348 6320 8406 6330
rect 8348 5934 8406 5948
rect 8684 6320 8742 6330
rect 8684 5934 8742 5948
rect 9020 6320 9078 6330
rect 11302 6324 11318 6614
rect 11542 6324 11560 6614
rect 17672 6614 17930 6630
rect 11302 6304 11560 6324
rect 13710 6320 13768 6330
rect 9020 5934 9078 5948
rect 13710 5934 13768 5948
rect 14046 6320 14104 6330
rect 14046 5934 14104 5948
rect 14382 6320 14440 6330
rect 14382 5934 14440 5948
rect 14718 6320 14776 6330
rect 14718 5934 14776 5948
rect 15054 6320 15112 6330
rect 15054 5934 15112 5948
rect 15390 6320 15448 6330
rect 17672 6324 17688 6614
rect 17912 6324 17930 6614
rect 24012 6614 24270 6630
rect 17672 6304 17930 6324
rect 20080 6320 20138 6330
rect 15390 5934 15448 5948
rect 20080 5934 20138 5948
rect 20416 6320 20474 6330
rect 20416 5934 20474 5948
rect 20752 6320 20810 6330
rect 20752 5934 20810 5948
rect 21088 6320 21146 6330
rect 21088 5934 21146 5948
rect 21424 6320 21482 6330
rect 21424 5934 21482 5948
rect 21760 6320 21818 6330
rect 24012 6324 24028 6614
rect 24252 6324 24270 6614
rect 29160 6486 31170 6670
rect 24012 6304 24270 6324
rect 29338 6320 29396 6330
rect 21760 5934 21818 5948
rect 29338 5934 29396 5948
rect 29674 6320 29732 6330
rect 29674 5934 29732 5948
rect 30010 6320 30068 6330
rect 30010 5934 30068 5948
rect 30346 6320 30404 6330
rect 30346 5934 30404 5948
rect 30682 6320 30740 6330
rect 30682 5934 30740 5948
rect 31018 6320 31076 6330
rect 31018 5934 31076 5948
rect -2748 5884 -2690 5898
rect -1684 5806 2900 5836
rect -5208 5756 -2498 5786
rect -5208 5704 -5200 5756
rect -2518 5704 -2498 5756
rect -1684 5754 -1656 5806
rect -1208 5754 796 5806
rect 2880 5754 2900 5806
rect -1684 5724 2900 5754
rect 4686 5806 9270 5836
rect 4686 5754 4714 5806
rect 5162 5754 7166 5806
rect 9250 5754 9270 5806
rect 4686 5724 9270 5754
rect 11056 5806 15640 5836
rect 11056 5754 11084 5806
rect 11532 5754 13536 5806
rect 15620 5754 15640 5806
rect 11056 5724 15640 5754
rect 17426 5806 22010 5836
rect 17426 5754 17454 5806
rect 17902 5754 19906 5806
rect 21990 5754 22010 5806
rect 17426 5724 22010 5754
rect 23766 5806 31268 5836
rect 23766 5754 23794 5806
rect 24242 5754 29164 5806
rect 31248 5754 31268 5806
rect 23766 5724 31268 5754
rect 35578 5778 35668 8436
rect 35892 5778 35980 8480
rect 35578 5736 35980 5778
rect -5208 5674 -2498 5704
rect 2980 5662 3092 5672
rect -2418 5612 -2306 5622
rect -2418 5444 -2390 5612
rect -2334 5444 -2306 5612
rect 2980 5494 3008 5662
rect 3064 5494 3092 5662
rect 2980 5484 3092 5494
rect 9350 5662 9462 5672
rect 9350 5494 9378 5662
rect 9434 5494 9462 5662
rect 9350 5484 9462 5494
rect 15720 5662 15832 5672
rect 15720 5494 15748 5662
rect 15804 5494 15832 5662
rect 15720 5484 15832 5494
rect 22090 5662 22202 5672
rect 22090 5494 22118 5662
rect 22174 5494 22202 5662
rect 22090 5484 22202 5494
rect 31348 5662 31460 5672
rect 31348 5494 31376 5662
rect 31432 5494 31460 5662
rect 31348 5484 31460 5494
rect -2418 5434 -2306 5444
<< via2 >>
rect -4918 8654 -4862 8822
rect 480 8704 536 8872
rect -4598 7372 -4540 8348
rect -4194 7372 -4136 8348
rect -3790 7372 -3732 8348
rect -3386 7372 -3328 8348
rect -2982 7372 -2924 8348
rect -2578 7372 -2520 8348
rect -5226 6326 -5002 6616
rect -4428 5898 -4370 6874
rect -4092 5898 -4034 6874
rect -3756 5898 -3698 6874
rect -3420 5898 -3362 6874
rect -3084 5898 -3026 6874
rect -2748 5898 -2690 6874
rect -2212 6722 -1994 8580
rect 6850 8704 6906 8872
rect 800 7422 858 8398
rect 1204 7422 1262 8398
rect 1608 7422 1666 8398
rect 2012 7422 2070 8398
rect 2416 7422 2474 8398
rect 2820 7422 2878 8398
rect -1640 6772 -646 6884
rect 3572 6728 3684 8580
rect 13220 8704 13276 8872
rect 7170 7422 7228 8398
rect 7574 7422 7632 8398
rect 7978 7422 8036 8398
rect 8382 7422 8440 8398
rect 8786 7422 8844 8398
rect 9190 7422 9248 8398
rect 4730 6772 5724 6884
rect 9942 6728 10054 8580
rect 19590 8704 19646 8872
rect 13540 7422 13598 8398
rect 13944 7422 14002 8398
rect 14348 7422 14406 8398
rect 14752 7422 14810 8398
rect 15156 7422 15214 8398
rect 15560 7422 15618 8398
rect 11100 6772 12094 6884
rect 16312 6728 16424 8580
rect 28848 8704 28904 8872
rect 19910 7422 19968 8398
rect 20314 7422 20372 8398
rect 20718 7422 20776 8398
rect 21122 7422 21180 8398
rect 21526 7422 21584 8398
rect 21930 7422 21988 8398
rect 17470 6772 18464 6884
rect 22682 6728 22794 8580
rect 29168 7422 29226 8398
rect 29572 7422 29630 8398
rect 29976 7422 30034 8398
rect 30380 7422 30438 8398
rect 30784 7422 30842 8398
rect 31188 7422 31246 8398
rect 23810 6772 24804 6884
rect -1422 6324 -1198 6614
rect 970 5948 1028 6320
rect 1306 5948 1364 6320
rect 1642 5948 1700 6320
rect 1978 5948 2036 6320
rect 2314 5948 2372 6320
rect 2650 5948 2708 6320
rect 4948 6324 5172 6614
rect 7340 5948 7398 6320
rect 7676 5948 7734 6320
rect 8012 5948 8070 6320
rect 8348 5948 8406 6320
rect 8684 5948 8742 6320
rect 9020 5948 9078 6320
rect 11318 6324 11542 6614
rect 13710 5948 13768 6320
rect 14046 5948 14104 6320
rect 14382 5948 14440 6320
rect 14718 5948 14776 6320
rect 15054 5948 15112 6320
rect 15390 5948 15448 6320
rect 17688 6324 17912 6614
rect 20080 5948 20138 6320
rect 20416 5948 20474 6320
rect 20752 5948 20810 6320
rect 21088 5948 21146 6320
rect 21424 5948 21482 6320
rect 21760 5948 21818 6320
rect 24028 6324 24252 6614
rect 29338 5948 29396 6320
rect 29674 5948 29732 6320
rect 30010 5948 30068 6320
rect 30346 5948 30404 6320
rect 30682 5948 30740 6320
rect 31018 5948 31076 6320
rect 35668 5778 35892 8480
rect -2390 5444 -2334 5612
rect 3008 5494 3064 5662
rect 9378 5494 9434 5662
rect 15748 5494 15804 5662
rect 22118 5494 22174 5662
rect 31376 5494 31432 5662
<< metal3 >>
rect -1584 8990 4496 15278
rect -1584 8926 -1556 8990
rect 4468 8926 4496 8990
rect -1584 8872 4496 8926
rect -5208 8822 -2000 8856
rect -5208 8776 -4918 8822
rect -4862 8776 -2000 8822
rect -5208 8706 -5202 8776
rect -2006 8706 -2000 8776
rect -5208 8654 -4918 8706
rect -4862 8700 -2000 8706
rect -1584 8704 480 8872
rect 536 8704 4496 8872
rect -4862 8654 -2302 8700
rect -1584 8676 4496 8704
rect 4786 8990 10866 15278
rect 4786 8926 4814 8990
rect 10838 8926 10866 8990
rect 4786 8872 10866 8926
rect 4786 8704 6850 8872
rect 6906 8704 10866 8872
rect 4786 8676 10866 8704
rect 11156 8990 17236 15278
rect 11156 8926 11184 8990
rect 17208 8926 17236 8990
rect 11156 8872 17236 8926
rect 11156 8704 13220 8872
rect 13276 8704 17236 8872
rect 11156 8676 17236 8704
rect 17526 8990 23606 15278
rect 17526 8926 17554 8990
rect 23578 8926 23606 8990
rect 17526 8872 23606 8926
rect 17526 8704 19590 8872
rect 19646 8704 23606 8872
rect 17526 8676 23606 8704
rect 23866 8990 29946 15278
rect 30186 9282 36266 15570
rect 30186 9218 30214 9282
rect 36238 9218 36266 9282
rect 30186 9198 36266 9218
rect 36346 15480 36586 15490
rect 36346 9580 36410 15480
rect 36522 9580 36586 15480
rect 23866 8926 23894 8990
rect 29918 8926 29946 8990
rect 23866 8906 29946 8926
rect 23866 8872 30848 8906
rect 23866 8704 28848 8872
rect 28904 8704 30848 8872
rect 23866 8676 30848 8704
rect -5208 8626 -2302 8654
rect -4604 8348 -4424 8626
rect -4604 7372 -4598 8348
rect -4540 7372 -4424 8348
rect -4604 6880 -4424 7372
rect -4200 8348 -4020 8360
rect -4200 7372 -4194 8348
rect -4136 7372 -4020 8348
rect -4604 6874 -4364 6880
rect -5242 6616 -4984 6632
rect -5242 6326 -5226 6616
rect -5002 6326 -4984 6616
rect -5242 6306 -4984 6326
rect -4604 5898 -4428 6874
rect -4370 5898 -4364 6874
rect -4604 5892 -4364 5898
rect -4200 6874 -4020 7372
rect -4200 5898 -4092 6874
rect -4034 5898 -4020 6874
rect -4200 5638 -4020 5898
rect -3796 8348 -3616 8626
rect -3796 7372 -3790 8348
rect -3732 7372 -3616 8348
rect -3796 6874 -3616 7372
rect -3796 5898 -3756 6874
rect -3698 5898 -3616 6874
rect -3796 5892 -3616 5898
rect -3442 8348 -3262 8360
rect -3442 7372 -3386 8348
rect -3328 7372 -3262 8348
rect -3442 6874 -3262 7372
rect -3442 5898 -3420 6874
rect -3362 5898 -3262 6874
rect -3442 5638 -3262 5898
rect -3098 8348 -2918 8626
rect -1684 8592 -604 8596
rect -2224 8580 -604 8592
rect -3098 7372 -2982 8348
rect -2924 7372 -2918 8348
rect -3098 6874 -2918 7372
rect -3098 5898 -3084 6874
rect -3026 5898 -2918 6874
rect -3098 5892 -2918 5898
rect -2754 8348 -2514 8360
rect -2754 7372 -2578 8348
rect -2520 7372 -2514 8348
rect -2754 7360 -2514 7372
rect -2754 6874 -2568 7360
rect -2754 5898 -2748 6874
rect -2690 5898 -2568 6874
rect -2224 6722 -2212 8580
rect -1994 6884 -604 8580
rect -1994 6772 -1640 6884
rect -646 6772 -604 6884
rect -1994 6722 -604 6772
rect -2224 6710 -604 6722
rect 794 8398 974 8676
rect 794 7422 800 8398
rect 858 7422 974 8398
rect 794 6930 974 7422
rect 1198 8398 1378 8410
rect 1198 7422 1204 8398
rect 1262 7422 1378 8398
rect -1438 6614 -1180 6630
rect -1438 6324 -1422 6614
rect -1198 6324 -1180 6614
rect -1438 6304 -1180 6324
rect 794 6320 1034 6930
rect 794 5948 970 6320
rect 1028 5948 1034 6320
rect 794 5942 1034 5948
rect 1198 6320 1378 7422
rect 1198 5948 1306 6320
rect 1364 5948 1378 6320
rect -2754 5638 -2568 5898
rect 1198 5688 1378 5948
rect 1602 8398 1782 8676
rect 1602 7422 1608 8398
rect 1666 7422 1782 8398
rect 1602 6320 1782 7422
rect 1602 5948 1642 6320
rect 1700 5948 1782 6320
rect 1602 5942 1782 5948
rect 1956 8398 2136 8410
rect 1956 7422 2012 8398
rect 2070 7422 2136 8398
rect 1956 6320 2136 7422
rect 1956 5948 1978 6320
rect 2036 5948 2136 6320
rect 1956 5688 2136 5948
rect 2300 8398 2480 8676
rect 3516 8580 5766 8596
rect 2300 7422 2416 8398
rect 2474 7422 2480 8398
rect 2300 6320 2480 7422
rect 2300 5948 2314 6320
rect 2372 5948 2480 6320
rect 2300 5942 2480 5948
rect 2644 8398 2884 8410
rect 2644 7422 2820 8398
rect 2878 7422 2884 8398
rect 2644 7410 2884 7422
rect 2644 6320 2830 7410
rect 3516 6728 3572 8580
rect 3684 6884 5766 8580
rect 3684 6772 4730 6884
rect 5724 6772 5766 6884
rect 3684 6728 5766 6772
rect 3516 6710 5766 6728
rect 7164 8398 7344 8676
rect 7164 7422 7170 8398
rect 7228 7422 7344 8398
rect 7164 6930 7344 7422
rect 7568 8398 7748 8410
rect 7568 7422 7574 8398
rect 7632 7422 7748 8398
rect 2644 5948 2650 6320
rect 2708 5948 2830 6320
rect 4932 6614 5190 6630
rect 4932 6324 4948 6614
rect 5172 6324 5190 6614
rect 4932 6304 5190 6324
rect 7164 6320 7404 6930
rect 2644 5688 2830 5948
rect 7164 5948 7340 6320
rect 7398 5948 7404 6320
rect 7164 5942 7404 5948
rect 7568 6320 7748 7422
rect 7568 5948 7676 6320
rect 7734 5948 7748 6320
rect 7568 5688 7748 5948
rect 7972 8398 8152 8676
rect 7972 7422 7978 8398
rect 8036 7422 8152 8398
rect 7972 6320 8152 7422
rect 7972 5948 8012 6320
rect 8070 5948 8152 6320
rect 7972 5942 8152 5948
rect 8326 8398 8506 8410
rect 8326 7422 8382 8398
rect 8440 7422 8506 8398
rect 8326 6320 8506 7422
rect 8326 5948 8348 6320
rect 8406 5948 8506 6320
rect 8326 5688 8506 5948
rect 8670 8398 8850 8676
rect 9886 8580 12136 8596
rect 8670 7422 8786 8398
rect 8844 7422 8850 8398
rect 8670 6320 8850 7422
rect 8670 5948 8684 6320
rect 8742 5948 8850 6320
rect 8670 5942 8850 5948
rect 9014 8398 9254 8410
rect 9014 7422 9190 8398
rect 9248 7422 9254 8398
rect 9014 7410 9254 7422
rect 9014 6320 9200 7410
rect 9886 6728 9942 8580
rect 10054 6884 12136 8580
rect 10054 6772 11100 6884
rect 12094 6772 12136 6884
rect 10054 6728 12136 6772
rect 9886 6710 12136 6728
rect 13534 8398 13714 8676
rect 13534 7422 13540 8398
rect 13598 7422 13714 8398
rect 13534 6930 13714 7422
rect 13938 8398 14118 8410
rect 13938 7422 13944 8398
rect 14002 7422 14118 8398
rect 9014 5948 9020 6320
rect 9078 5948 9200 6320
rect 11302 6614 11560 6630
rect 11302 6324 11318 6614
rect 11542 6324 11560 6614
rect 11302 6304 11560 6324
rect 13534 6320 13774 6930
rect 9014 5688 9200 5948
rect 13534 5948 13710 6320
rect 13768 5948 13774 6320
rect 13534 5942 13774 5948
rect 13938 6320 14118 7422
rect 13938 5948 14046 6320
rect 14104 5948 14118 6320
rect 13938 5688 14118 5948
rect 14342 8398 14522 8676
rect 14342 7422 14348 8398
rect 14406 7422 14522 8398
rect 14342 6320 14522 7422
rect 14342 5948 14382 6320
rect 14440 5948 14522 6320
rect 14342 5942 14522 5948
rect 14696 8398 14876 8410
rect 14696 7422 14752 8398
rect 14810 7422 14876 8398
rect 14696 6320 14876 7422
rect 14696 5948 14718 6320
rect 14776 5948 14876 6320
rect 14696 5688 14876 5948
rect 15040 8398 15220 8676
rect 16256 8580 18506 8596
rect 15040 7422 15156 8398
rect 15214 7422 15220 8398
rect 15040 6320 15220 7422
rect 15040 5948 15054 6320
rect 15112 5948 15220 6320
rect 15040 5942 15220 5948
rect 15384 8398 15624 8410
rect 15384 7422 15560 8398
rect 15618 7422 15624 8398
rect 15384 7410 15624 7422
rect 15384 6320 15570 7410
rect 16256 6728 16312 8580
rect 16424 6884 18506 8580
rect 16424 6772 17470 6884
rect 18464 6772 18506 6884
rect 16424 6728 18506 6772
rect 16256 6710 18506 6728
rect 19904 8398 20084 8676
rect 19904 7422 19910 8398
rect 19968 7422 20084 8398
rect 19904 6930 20084 7422
rect 20308 8398 20488 8410
rect 20308 7422 20314 8398
rect 20372 7422 20488 8398
rect 15384 5948 15390 6320
rect 15448 5948 15570 6320
rect 17672 6614 17930 6630
rect 17672 6324 17688 6614
rect 17912 6324 17930 6614
rect 17672 6304 17930 6324
rect 19904 6320 20144 6930
rect 15384 5688 15570 5948
rect 19904 5948 20080 6320
rect 20138 5948 20144 6320
rect 19904 5942 20144 5948
rect 20308 6320 20488 7422
rect 20308 5948 20416 6320
rect 20474 5948 20488 6320
rect 20308 5688 20488 5948
rect 20712 8398 20892 8676
rect 20712 7422 20718 8398
rect 20776 7422 20892 8398
rect 20712 6320 20892 7422
rect 20712 5948 20752 6320
rect 20810 5948 20892 6320
rect 20712 5942 20892 5948
rect 21066 8398 21246 8410
rect 21066 7422 21122 8398
rect 21180 7422 21246 8398
rect 21066 6320 21246 7422
rect 21066 5948 21088 6320
rect 21146 5948 21246 6320
rect 21066 5688 21246 5948
rect 21410 8398 21590 8676
rect 22626 8580 24846 8596
rect 21410 7422 21526 8398
rect 21584 7422 21590 8398
rect 21410 6320 21590 7422
rect 21410 5948 21424 6320
rect 21482 5948 21590 6320
rect 21410 5942 21590 5948
rect 21754 8398 21994 8410
rect 21754 7422 21930 8398
rect 21988 7422 21994 8398
rect 21754 7410 21994 7422
rect 21754 6320 21940 7410
rect 22626 6728 22682 8580
rect 22794 6884 24846 8580
rect 22794 6772 23810 6884
rect 24804 6772 24846 6884
rect 22794 6728 24846 6772
rect 22626 6710 24846 6728
rect 29162 8398 29342 8676
rect 29162 7422 29168 8398
rect 29226 7422 29342 8398
rect 29162 6930 29342 7422
rect 29566 8398 29746 8410
rect 29566 7422 29572 8398
rect 29630 7422 29746 8398
rect 21754 5948 21760 6320
rect 21818 5948 21940 6320
rect 24012 6614 24270 6630
rect 24012 6324 24028 6614
rect 24252 6324 24270 6614
rect 24012 6304 24270 6324
rect 29162 6320 29402 6930
rect 21754 5688 21940 5948
rect 29162 5948 29338 6320
rect 29396 5948 29402 6320
rect 29162 5942 29402 5948
rect 29566 6320 29746 7422
rect 29566 5948 29674 6320
rect 29732 5948 29746 6320
rect 29566 5688 29746 5948
rect 29970 8398 30150 8676
rect 29970 7422 29976 8398
rect 30034 7422 30150 8398
rect 29970 6320 30150 7422
rect 29970 5948 30010 6320
rect 30068 5948 30150 6320
rect 29970 5942 30150 5948
rect 30324 8398 30504 8410
rect 30324 7422 30380 8398
rect 30438 7422 30504 8398
rect 30324 6320 30504 7422
rect 30324 5948 30346 6320
rect 30404 5948 30504 6320
rect 30324 5688 30504 5948
rect 30668 8398 30848 8676
rect 36346 8536 36586 9580
rect 35578 8480 36658 8536
rect 30668 7422 30784 8398
rect 30842 7422 30848 8398
rect 30668 6320 30848 7422
rect 30668 5948 30682 6320
rect 30740 5948 30848 6320
rect 30668 5942 30848 5948
rect 31012 8398 31252 8410
rect 31012 7422 31188 8398
rect 31246 7422 31252 8398
rect 31012 7410 31252 7422
rect 31012 6320 31198 7410
rect 31012 5948 31018 6320
rect 31076 5948 31198 6320
rect 31012 5688 31198 5948
rect 35578 5778 35668 8480
rect 35892 5778 36658 8480
rect 35578 5736 36658 5778
rect -1584 5662 4496 5688
rect -5208 5612 -2000 5638
rect -5208 5554 -2390 5612
rect -2334 5554 -2000 5612
rect -5208 5484 -5202 5554
rect -2006 5484 -2000 5554
rect -5208 5444 -2390 5484
rect -2334 5444 -2000 5484
rect -1584 5604 3008 5662
rect 3064 5604 4496 5662
rect -1584 5534 -1578 5604
rect 4486 5534 4496 5604
rect -1584 5494 3008 5534
rect 3064 5494 4496 5534
rect -1584 5448 4496 5494
rect 4786 5662 10866 5688
rect 4786 5604 9378 5662
rect 9434 5604 10866 5662
rect 4786 5534 4792 5604
rect 10856 5534 10866 5604
rect 4786 5494 9378 5534
rect 9434 5494 10866 5534
rect 4786 5448 10866 5494
rect 11156 5662 17236 5688
rect 11156 5604 15748 5662
rect 15804 5604 17236 5662
rect 11156 5534 11162 5604
rect 17226 5534 17236 5604
rect 11156 5494 15748 5534
rect 15804 5494 17236 5534
rect 11156 5448 17236 5494
rect 17526 5662 23606 5688
rect 17526 5604 22118 5662
rect 22174 5604 23606 5662
rect 17526 5534 17532 5604
rect 23596 5534 23606 5604
rect 17526 5494 22118 5534
rect 22174 5494 23606 5534
rect 17526 5448 23606 5494
rect 23866 5662 31476 5688
rect 23866 5604 31376 5662
rect 31432 5604 31476 5662
rect 23866 5534 23872 5604
rect 31470 5534 31476 5604
rect 23866 5494 31376 5534
rect 31432 5494 31476 5534
rect 23866 5448 31476 5494
rect -5208 5432 -2000 5444
rect -1584 -920 4496 5368
rect -1584 -984 -1556 -920
rect 4468 -984 4496 -920
rect -1584 -1004 4496 -984
rect 4786 -920 10866 5368
rect 4786 -984 4814 -920
rect 10838 -984 10866 -920
rect 4786 -1004 10866 -984
rect 11156 -920 17236 5368
rect 11156 -984 11184 -920
rect 17208 -984 17236 -920
rect 11156 -1004 17236 -984
rect 17526 -920 23606 5368
rect 17526 -984 17554 -920
rect 23578 -984 23606 -920
rect 17526 -1004 23606 -984
rect 23866 -920 29946 5368
rect 23866 -984 23894 -920
rect 29918 -984 29946 -920
rect 23866 -1004 29946 -984
rect 30186 5348 36266 5368
rect 30186 5284 30214 5348
rect 36238 5284 36266 5348
rect 30186 -1004 36266 5284
rect 36346 4986 36586 5736
rect 36346 -914 36410 4986
rect 36522 -914 36586 4986
rect 36346 -1004 36586 -914
<< via3 >>
rect -1556 8926 4468 8990
rect -5202 8706 -4918 8776
rect -4918 8706 -4862 8776
rect -4862 8706 -2006 8776
rect 4814 8926 10838 8990
rect 11184 8926 17208 8990
rect 17554 8926 23578 8990
rect 30214 9218 36238 9282
rect 36410 9580 36522 15480
rect 23894 8926 29918 8990
rect -5226 6326 -5002 6616
rect -1422 6324 -1198 6614
rect 4948 6324 5172 6614
rect 11318 6324 11542 6614
rect 17688 6324 17912 6614
rect 24028 6324 24252 6614
rect -5202 5484 -2390 5554
rect -2390 5484 -2334 5554
rect -2334 5484 -2006 5554
rect -1578 5534 3008 5604
rect 3008 5534 3064 5604
rect 3064 5534 4486 5604
rect 4792 5534 9378 5604
rect 9378 5534 9434 5604
rect 9434 5534 10856 5604
rect 11162 5534 15748 5604
rect 15748 5534 15804 5604
rect 15804 5534 17226 5604
rect 17532 5534 22118 5604
rect 22118 5534 22174 5604
rect 22174 5534 23596 5604
rect 23872 5534 31376 5604
rect 31376 5534 31432 5604
rect 31432 5534 31470 5604
rect -1556 -984 4468 -920
rect 4814 -984 10838 -920
rect 11184 -984 17208 -920
rect 17554 -984 23578 -920
rect 23894 -984 29918 -920
rect 30214 5284 36238 5348
rect 36410 -914 36522 4986
<< mimcap >>
rect 30226 15490 36226 15530
rect -1544 15198 4456 15238
rect -1544 9278 -1504 15198
rect 4416 9278 4456 15198
rect -1544 9238 4456 9278
rect 4826 15198 10826 15238
rect 4826 9278 4866 15198
rect 10786 9278 10826 15198
rect 4826 9238 10826 9278
rect 11196 15198 17196 15238
rect 11196 9278 11236 15198
rect 17156 9278 17196 15198
rect 11196 9238 17196 9278
rect 17566 15198 23566 15238
rect 17566 9278 17606 15198
rect 23526 9278 23566 15198
rect 17566 9238 23566 9278
rect 23906 15198 29906 15238
rect 23906 9278 23946 15198
rect 29866 9278 29906 15198
rect 30226 9570 30266 15490
rect 36186 9570 36226 15490
rect 30226 9530 36226 9570
rect 23906 9238 29906 9278
rect -1544 5288 4456 5328
rect -1544 -632 -1504 5288
rect 4416 -632 4456 5288
rect -1544 -672 4456 -632
rect 4826 5288 10826 5328
rect 4826 -632 4866 5288
rect 10786 -632 10826 5288
rect 4826 -672 10826 -632
rect 11196 5288 17196 5328
rect 11196 -632 11236 5288
rect 17156 -632 17196 5288
rect 11196 -672 17196 -632
rect 17566 5288 23566 5328
rect 17566 -632 17606 5288
rect 23526 -632 23566 5288
rect 17566 -672 23566 -632
rect 23906 5288 29906 5328
rect 23906 -632 23946 5288
rect 29866 -632 29906 5288
rect 23906 -672 29906 -632
rect 30226 4996 36226 5036
rect 30226 -924 30266 4996
rect 36186 -924 36226 4996
rect 30226 -964 36226 -924
<< mimcapcontact >>
rect -1504 9278 4416 15198
rect 4866 9278 10786 15198
rect 11236 9278 17156 15198
rect 17606 9278 23526 15198
rect 23946 9278 29866 15198
rect 30266 9570 36186 15490
rect -1504 -632 4416 5288
rect 4866 -632 10786 5288
rect 11236 -632 17156 5288
rect 17606 -632 23526 5288
rect 23946 -632 29866 5288
rect 30266 -924 36186 4996
<< metal4 >>
rect -5208 15298 29866 16378
rect -5208 8776 -2000 15298
rect -1504 15199 4416 15298
rect 4866 15199 10786 15298
rect 11236 15199 17156 15298
rect 17606 15199 23526 15298
rect 23946 15199 29866 15298
rect 30265 15490 36187 15491
rect -1505 15198 4417 15199
rect -1505 9278 -1504 15198
rect 4416 9278 4417 15198
rect -1505 9277 4417 9278
rect 4865 15198 10787 15199
rect 4865 9278 4866 15198
rect 10786 9278 10787 15198
rect 4865 9277 10787 9278
rect 11235 15198 17157 15199
rect 11235 9278 11236 15198
rect 17156 9278 17157 15198
rect 11235 9277 17157 9278
rect 17605 15198 23527 15199
rect 17605 9278 17606 15198
rect 23526 9278 23527 15198
rect 17605 9277 23527 9278
rect 23945 15198 29867 15199
rect 23945 9278 23946 15198
rect 29866 9278 29867 15198
rect 30265 9570 30266 15490
rect 36186 15480 36528 15490
rect 36186 9580 36410 15480
rect 36522 9580 36528 15480
rect 36186 9570 36528 9580
rect 30265 9569 36187 9570
rect 23945 9277 29867 9278
rect 30198 9282 36254 9298
rect 30198 9218 30214 9282
rect 36238 9218 36254 9282
rect 30198 9202 36254 9218
rect -1572 8990 4484 9006
rect -1572 8926 -1556 8990
rect 4468 8926 4484 8990
rect -1572 8910 4484 8926
rect 4798 8990 10854 9006
rect 4798 8926 4814 8990
rect 10838 8926 10854 8990
rect 4798 8910 10854 8926
rect 11168 8990 17224 9006
rect 11168 8926 11184 8990
rect 17208 8926 17224 8990
rect 11168 8910 17224 8926
rect 17538 8990 23594 9006
rect 17538 8926 17554 8990
rect 23578 8926 23594 8990
rect 17538 8910 23594 8926
rect 23878 8990 29934 9006
rect 23878 8926 23894 8990
rect 29918 8926 29934 8990
rect 23878 8910 29934 8926
rect -5208 8706 -5202 8776
rect -2006 8706 -2000 8776
rect -5208 8700 -2000 8706
rect -5242 6664 -4984 6666
rect 33010 6664 33370 9202
rect -5242 6616 33370 6664
rect -5242 6326 -5226 6616
rect -5002 6614 33370 6616
rect -5002 6326 -1422 6614
rect -5242 6324 -1422 6326
rect -1198 6324 4948 6614
rect 5172 6324 11318 6614
rect 11542 6324 17688 6614
rect 17912 6324 24028 6614
rect 24252 6324 33370 6614
rect -5242 6306 33370 6324
rect -1438 6304 -1180 6306
rect 4932 6304 5190 6306
rect 11302 6304 11560 6306
rect 17672 6304 17930 6306
rect 24012 6304 33370 6306
rect -1584 5604 4496 5610
rect -5208 5554 -2000 5560
rect -5208 5484 -5202 5554
rect -2006 5484 -2000 5554
rect -5208 -1024 -2000 5484
rect -1584 5534 -1578 5604
rect 4486 5534 4496 5604
rect -1584 5288 4496 5534
rect -1584 5284 -1504 5288
rect -1505 -632 -1504 5284
rect 4416 5284 4496 5288
rect 4786 5604 10866 5610
rect 4786 5534 4792 5604
rect 10856 5534 10866 5604
rect 4786 5288 10866 5534
rect 4786 5284 4866 5288
rect 4416 -632 4417 5284
rect -1505 -633 4417 -632
rect 4865 -632 4866 5284
rect 10786 5284 10866 5288
rect 11156 5604 17236 5610
rect 11156 5534 11162 5604
rect 17226 5534 17236 5604
rect 11156 5288 17236 5534
rect 11156 5284 11236 5288
rect 10786 -632 10787 5284
rect 4865 -633 10787 -632
rect 11235 -632 11236 5284
rect 17156 5284 17236 5288
rect 17526 5604 23606 5610
rect 17526 5534 17532 5604
rect 23596 5534 23606 5604
rect 17526 5288 23606 5534
rect 17526 5284 17606 5288
rect 17156 -632 17157 5284
rect 11235 -633 17157 -632
rect 17605 -632 17606 5284
rect 23526 5284 23606 5288
rect 23866 5604 31476 5610
rect 23866 5534 23872 5604
rect 31470 5534 31476 5604
rect 23866 5428 31476 5534
rect 23866 5288 29946 5428
rect 33010 5364 33370 6304
rect 23866 5284 23946 5288
rect 23526 -632 23527 5284
rect 17605 -633 23527 -632
rect 23945 -632 23946 5284
rect 29866 5284 29946 5288
rect 30198 5348 36254 5364
rect 30198 5284 30214 5348
rect 36238 5284 36254 5348
rect 29866 -632 29867 5284
rect 30198 5268 36254 5284
rect 23945 -633 29867 -632
rect 30265 4996 36187 4997
rect -1572 -910 4484 -904
rect 4798 -910 10854 -904
rect 11168 -910 17224 -904
rect 17538 -910 23594 -904
rect -1684 -920 4598 -910
rect -1684 -984 -1556 -920
rect 4468 -984 4598 -920
rect -1684 -1024 4598 -984
rect 4686 -920 10968 -910
rect 4686 -984 4814 -920
rect 10838 -984 10968 -920
rect 4686 -1024 10968 -984
rect 11056 -920 17338 -910
rect 11056 -984 11184 -920
rect 17208 -984 17338 -920
rect 11056 -1024 17338 -984
rect 17426 -920 23708 -910
rect 17426 -984 17554 -920
rect 23578 -984 23708 -920
rect 17426 -1000 23708 -984
rect 23878 -920 29934 -904
rect 23878 -984 23894 -920
rect 29918 -984 29934 -920
rect 30265 -924 30266 4996
rect 36186 4986 36528 4996
rect 36186 -914 36410 4986
rect 36522 -914 36528 4986
rect 36186 -924 36528 -914
rect 30265 -925 36187 -924
rect 23878 -1000 29934 -984
rect 17426 -1024 29866 -1000
rect -5208 -2104 29866 -1024
<< labels >>
flabel metal4 -5208 15302 29866 16378 0 FreeMono 4800 0 0 0 vinp
port 1 nsew
flabel metal4 -5208 -2104 29866 -1024 0 FreeMono 4800 0 0 0 vinn
port 2 nsew
flabel metal1 -5242 5674 -4984 8522 0 FreeMono 1600 90 0 0 vss
port 0 nsew
flabel metal3 35578 5736 36658 8536 0 FreeMono 1920 0 0 0 vrec
port 3 nsew
<< end >>
