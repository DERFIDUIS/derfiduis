magic
tech sky130A
magscale 1 2
timestamp 1680254065
<< nwell >>
rect -633 -591 633 591
<< varactor >>
rect -500 -500 500 500
<< nsubdiff >>
rect -597 476 -500 500
rect -597 -476 -585 476
rect -551 -476 -500 476
rect -597 -500 -500 -476
rect 500 476 597 500
rect 500 -476 551 476
rect 585 -476 597 476
rect 500 -500 597 -476
<< nsubdiffcont >>
rect -585 -476 -551 476
rect 551 -476 585 476
<< poly >>
rect -500 572 500 588
rect -500 538 -484 572
rect 484 538 500 572
rect -500 500 500 538
rect -500 -538 500 -500
rect -500 -572 -484 -538
rect 484 -572 500 -538
rect -500 -588 500 -572
<< polycont >>
rect -484 538 484 572
rect -484 -572 484 -538
<< locali >>
rect -500 538 -484 572
rect 484 538 500 572
rect -585 476 -551 492
rect -585 -492 -551 -476
rect 551 476 585 492
rect 551 -492 585 -476
rect -500 -572 -484 -538
rect 484 -572 500 -538
<< viali >>
rect -484 538 484 572
rect -585 -476 -551 476
rect 551 -476 585 476
rect -484 -572 484 -538
<< metal1 >>
rect -496 572 496 578
rect -496 538 -484 572
rect 484 538 496 572
rect -496 532 496 538
rect -591 476 -545 488
rect -591 -476 -585 476
rect -551 -476 -545 476
rect -591 -488 -545 -476
rect 545 476 591 488
rect 545 -476 551 476
rect 585 -476 591 476
rect 545 -488 591 -476
rect -496 -538 496 -532
rect -496 -572 -484 -538
rect 484 -572 496 -538
rect -496 -578 496 -572
<< properties >>
string gencell sky130_fd_pr__cap_var_lvt
string library sky130
string parameters w 5.0 l 5.0 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.18 wmin 1.0 compatible {sky130_fd_pr__cap_var_lvt  sky130_fd_pr__cap_var_hvt sky130_fd_pr__cap_var} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
